magic
tech sky130A
timestamp 1723858470
<< properties >>
string GDS_END 6518
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 6130
<< end >>

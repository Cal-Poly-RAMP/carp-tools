magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< metal2 >>
rect 356 51378 412 51387
rect 356 51313 412 51322
rect 0 51199 28 51247
rect 356 51141 412 51150
rect 356 51076 412 51085
rect 0 50979 28 51027
rect 0 50883 28 50931
rect 356 50825 412 50834
rect 356 50760 412 50769
rect 0 50663 28 50711
rect 356 50588 412 50597
rect 356 50523 412 50532
rect 0 50409 28 50457
rect 356 50351 412 50360
rect 356 50286 412 50295
rect 0 50189 28 50237
rect 0 50093 28 50141
rect 356 50035 412 50044
rect 356 49970 412 49979
rect 0 49873 28 49921
rect 356 49798 412 49807
rect 356 49733 412 49742
rect 0 49619 28 49667
rect 356 49561 412 49570
rect 356 49496 412 49505
rect 0 49399 28 49447
rect 0 49303 28 49351
rect 356 49245 412 49254
rect 356 49180 412 49189
rect 0 49083 28 49131
rect 356 49008 412 49017
rect 356 48943 412 48952
rect 0 48829 28 48877
rect 356 48771 412 48780
rect 356 48706 412 48715
rect 0 48609 28 48657
rect 0 48513 28 48561
rect 356 48455 412 48464
rect 356 48390 412 48399
rect 0 48293 28 48341
rect 356 48218 412 48227
rect 356 48153 412 48162
rect 0 48039 28 48087
rect 356 47981 412 47990
rect 356 47916 412 47925
rect 0 47819 28 47867
rect 0 47723 28 47771
rect 356 47665 412 47674
rect 356 47600 412 47609
rect 0 47503 28 47551
rect 356 47428 412 47437
rect 356 47363 412 47372
rect 0 47249 28 47297
rect 356 47191 412 47200
rect 356 47126 412 47135
rect 0 47029 28 47077
rect 0 46933 28 46981
rect 356 46875 412 46884
rect 356 46810 412 46819
rect 0 46713 28 46761
rect 356 46638 412 46647
rect 356 46573 412 46582
rect 0 46459 28 46507
rect 356 46401 412 46410
rect 356 46336 412 46345
rect 0 46239 28 46287
rect 0 46143 28 46191
rect 356 46085 412 46094
rect 356 46020 412 46029
rect 0 45923 28 45971
rect 356 45848 412 45857
rect 356 45783 412 45792
rect 0 45669 28 45717
rect 356 45611 412 45620
rect 356 45546 412 45555
rect 0 45449 28 45497
rect 0 45353 28 45401
rect 356 45295 412 45304
rect 356 45230 412 45239
rect 0 45133 28 45181
rect 356 45058 412 45067
rect 356 44993 412 45002
rect 0 44879 28 44927
rect 356 44821 412 44830
rect 356 44756 412 44765
rect 0 44659 28 44707
rect 0 44563 28 44611
rect 356 44505 412 44514
rect 356 44440 412 44449
rect 0 44343 28 44391
rect 356 44268 412 44277
rect 356 44203 412 44212
rect 0 44089 28 44137
rect 356 44031 412 44040
rect 356 43966 412 43975
rect 0 43869 28 43917
rect 0 43773 28 43821
rect 356 43715 412 43724
rect 356 43650 412 43659
rect 0 43553 28 43601
rect 356 43478 412 43487
rect 356 43413 412 43422
rect 0 43299 28 43347
rect 356 43241 412 43250
rect 356 43176 412 43185
rect 0 43079 28 43127
rect 0 42983 28 43031
rect 356 42925 412 42934
rect 356 42860 412 42869
rect 0 42763 28 42811
rect 356 42688 412 42697
rect 356 42623 412 42632
rect 0 42509 28 42557
rect 356 42451 412 42460
rect 356 42386 412 42395
rect 0 42289 28 42337
rect 0 42193 28 42241
rect 356 42135 412 42144
rect 356 42070 412 42079
rect 0 41973 28 42021
rect 356 41898 412 41907
rect 356 41833 412 41842
rect 0 41719 28 41767
rect 356 41661 412 41670
rect 356 41596 412 41605
rect 0 41499 28 41547
rect 0 41403 28 41451
rect 356 41345 412 41354
rect 356 41280 412 41289
rect 0 41183 28 41231
rect 356 41108 412 41117
rect 356 41043 412 41052
rect 0 40929 28 40977
rect 356 40871 412 40880
rect 356 40806 412 40815
rect 0 40709 28 40757
rect 0 40613 28 40661
rect 356 40555 412 40564
rect 356 40490 412 40499
rect 0 40393 28 40441
rect 356 40318 412 40327
rect 356 40253 412 40262
rect 0 40139 28 40187
rect 356 40081 412 40090
rect 356 40016 412 40025
rect 0 39919 28 39967
rect 0 39823 28 39871
rect 356 39765 412 39774
rect 356 39700 412 39709
rect 0 39603 28 39651
rect 356 39528 412 39537
rect 356 39463 412 39472
rect 0 39349 28 39397
rect 356 39291 412 39300
rect 356 39226 412 39235
rect 0 39129 28 39177
rect 0 39033 28 39081
rect 356 38975 412 38984
rect 356 38910 412 38919
rect 0 38813 28 38861
rect 356 38738 412 38747
rect 356 38673 412 38682
rect 0 38559 28 38607
rect 356 38501 412 38510
rect 356 38436 412 38445
rect 0 38339 28 38387
rect 0 38243 28 38291
rect 356 38185 412 38194
rect 356 38120 412 38129
rect 0 38023 28 38071
rect 356 37948 412 37957
rect 356 37883 412 37892
rect 0 37769 28 37817
rect 356 37711 412 37720
rect 356 37646 412 37655
rect 0 37549 28 37597
rect 0 37453 28 37501
rect 356 37395 412 37404
rect 356 37330 412 37339
rect 0 37233 28 37281
rect 356 37158 412 37167
rect 356 37093 412 37102
rect 0 36979 28 37027
rect 356 36921 412 36930
rect 356 36856 412 36865
rect 0 36759 28 36807
rect 0 36663 28 36711
rect 356 36605 412 36614
rect 356 36540 412 36549
rect 0 36443 28 36491
rect 356 36368 412 36377
rect 356 36303 412 36312
rect 0 36189 28 36237
rect 356 36131 412 36140
rect 356 36066 412 36075
rect 0 35969 28 36017
rect 0 35873 28 35921
rect 356 35815 412 35824
rect 356 35750 412 35759
rect 0 35653 28 35701
rect 356 35578 412 35587
rect 356 35513 412 35522
rect 0 35399 28 35447
rect 356 35341 412 35350
rect 356 35276 412 35285
rect 0 35179 28 35227
rect 0 35083 28 35131
rect 356 35025 412 35034
rect 356 34960 412 34969
rect 0 34863 28 34911
rect 356 34788 412 34797
rect 356 34723 412 34732
rect 0 34609 28 34657
rect 356 34551 412 34560
rect 356 34486 412 34495
rect 0 34389 28 34437
rect 0 34293 28 34341
rect 356 34235 412 34244
rect 356 34170 412 34179
rect 0 34073 28 34121
rect 356 33998 412 34007
rect 356 33933 412 33942
rect 0 33819 28 33867
rect 356 33761 412 33770
rect 356 33696 412 33705
rect 0 33599 28 33647
rect 0 33503 28 33551
rect 356 33445 412 33454
rect 356 33380 412 33389
rect 0 33283 28 33331
rect 356 33208 412 33217
rect 356 33143 412 33152
rect 0 33029 28 33077
rect 356 32971 412 32980
rect 356 32906 412 32915
rect 0 32809 28 32857
rect 0 32713 28 32761
rect 356 32655 412 32664
rect 356 32590 412 32599
rect 0 32493 28 32541
rect 356 32418 412 32427
rect 356 32353 412 32362
rect 0 32239 28 32287
rect 356 32181 412 32190
rect 356 32116 412 32125
rect 0 32019 28 32067
rect 0 31923 28 31971
rect 356 31865 412 31874
rect 356 31800 412 31809
rect 0 31703 28 31751
rect 356 31628 412 31637
rect 356 31563 412 31572
rect 0 31449 28 31497
rect 356 31391 412 31400
rect 356 31326 412 31335
rect 0 31229 28 31277
rect 0 31133 28 31181
rect 356 31075 412 31084
rect 356 31010 412 31019
rect 0 30913 28 30961
rect 356 30838 412 30847
rect 356 30773 412 30782
rect 0 30659 28 30707
rect 356 30601 412 30610
rect 356 30536 412 30545
rect 0 30439 28 30487
rect 0 30343 28 30391
rect 356 30285 412 30294
rect 356 30220 412 30229
rect 0 30123 28 30171
rect 356 30048 412 30057
rect 356 29983 412 29992
rect 0 29869 28 29917
rect 356 29811 412 29820
rect 356 29746 412 29755
rect 0 29649 28 29697
rect 0 29553 28 29601
rect 356 29495 412 29504
rect 356 29430 412 29439
rect 0 29333 28 29381
rect 356 29258 412 29267
rect 356 29193 412 29202
rect 0 29079 28 29127
rect 356 29021 412 29030
rect 356 28956 412 28965
rect 0 28859 28 28907
rect 0 28763 28 28811
rect 356 28705 412 28714
rect 356 28640 412 28649
rect 0 28543 28 28591
rect 356 28468 412 28477
rect 356 28403 412 28412
rect 0 28289 28 28337
rect 356 28231 412 28240
rect 356 28166 412 28175
rect 0 28069 28 28117
rect 0 27973 28 28021
rect 356 27915 412 27924
rect 356 27850 412 27859
rect 0 27753 28 27801
rect 356 27678 412 27687
rect 356 27613 412 27622
rect 0 27499 28 27547
rect 356 27441 412 27450
rect 356 27376 412 27385
rect 0 27279 28 27327
rect 0 27183 28 27231
rect 356 27125 412 27134
rect 356 27060 412 27069
rect 0 26963 28 27011
rect 356 26888 412 26897
rect 356 26823 412 26832
rect 0 26709 28 26757
rect 356 26651 412 26660
rect 356 26586 412 26595
rect 0 26489 28 26537
rect 0 26393 28 26441
rect 356 26335 412 26344
rect 356 26270 412 26279
rect 0 26173 28 26221
rect 356 26098 412 26107
rect 356 26033 412 26042
rect 0 25919 28 25967
rect 356 25861 412 25870
rect 356 25796 412 25805
rect 0 25699 28 25747
rect 0 25603 28 25651
rect 356 25545 412 25554
rect 356 25480 412 25489
rect 0 25383 28 25431
rect 356 25308 412 25317
rect 356 25243 412 25252
rect 0 25129 28 25177
rect 356 25071 412 25080
rect 356 25006 412 25015
rect 0 24909 28 24957
rect 0 24813 28 24861
rect 356 24755 412 24764
rect 356 24690 412 24699
rect 0 24593 28 24641
rect 356 24518 412 24527
rect 356 24453 412 24462
rect 0 24339 28 24387
rect 356 24281 412 24290
rect 356 24216 412 24225
rect 0 24119 28 24167
rect 0 24023 28 24071
rect 356 23965 412 23974
rect 356 23900 412 23909
rect 0 23803 28 23851
rect 356 23728 412 23737
rect 356 23663 412 23672
rect 0 23549 28 23597
rect 356 23491 412 23500
rect 356 23426 412 23435
rect 0 23329 28 23377
rect 0 23233 28 23281
rect 356 23175 412 23184
rect 356 23110 412 23119
rect 0 23013 28 23061
rect 356 22938 412 22947
rect 356 22873 412 22882
rect 0 22759 28 22807
rect 356 22701 412 22710
rect 356 22636 412 22645
rect 0 22539 28 22587
rect 0 22443 28 22491
rect 356 22385 412 22394
rect 356 22320 412 22329
rect 0 22223 28 22271
rect 356 22148 412 22157
rect 356 22083 412 22092
rect 0 21969 28 22017
rect 356 21911 412 21920
rect 356 21846 412 21855
rect 0 21749 28 21797
rect 0 21653 28 21701
rect 356 21595 412 21604
rect 356 21530 412 21539
rect 0 21433 28 21481
rect 356 21358 412 21367
rect 356 21293 412 21302
rect 0 21179 28 21227
rect 356 21121 412 21130
rect 356 21056 412 21065
rect 0 20959 28 21007
rect 0 20863 28 20911
rect 356 20805 412 20814
rect 356 20740 412 20749
rect 0 20643 28 20691
rect 356 20568 412 20577
rect 356 20503 412 20512
rect 0 20389 28 20437
rect 356 20331 412 20340
rect 356 20266 412 20275
rect 0 20169 28 20217
rect 0 20073 28 20121
rect 356 20015 412 20024
rect 356 19950 412 19959
rect 0 19853 28 19901
rect 356 19778 412 19787
rect 356 19713 412 19722
rect 0 19599 28 19647
rect 356 19541 412 19550
rect 356 19476 412 19485
rect 0 19379 28 19427
rect 0 19283 28 19331
rect 356 19225 412 19234
rect 356 19160 412 19169
rect 0 19063 28 19111
rect 356 18988 412 18997
rect 356 18923 412 18932
rect 0 18809 28 18857
rect 356 18751 412 18760
rect 356 18686 412 18695
rect 0 18589 28 18637
rect 0 18493 28 18541
rect 356 18435 412 18444
rect 356 18370 412 18379
rect 0 18273 28 18321
rect 356 18198 412 18207
rect 356 18133 412 18142
rect 0 18019 28 18067
rect 356 17961 412 17970
rect 356 17896 412 17905
rect 0 17799 28 17847
rect 0 17703 28 17751
rect 356 17645 412 17654
rect 356 17580 412 17589
rect 0 17483 28 17531
rect 356 17408 412 17417
rect 356 17343 412 17352
rect 0 17229 28 17277
rect 356 17171 412 17180
rect 356 17106 412 17115
rect 0 17009 28 17057
rect 0 16913 28 16961
rect 356 16855 412 16864
rect 356 16790 412 16799
rect 0 16693 28 16741
rect 356 16618 412 16627
rect 356 16553 412 16562
rect 0 16439 28 16487
rect 356 16381 412 16390
rect 356 16316 412 16325
rect 0 16219 28 16267
rect 0 16123 28 16171
rect 356 16065 412 16074
rect 356 16000 412 16009
rect 0 15903 28 15951
rect 356 15828 412 15837
rect 356 15763 412 15772
rect 0 15649 28 15697
rect 356 15591 412 15600
rect 356 15526 412 15535
rect 0 15429 28 15477
rect 0 15333 28 15381
rect 356 15275 412 15284
rect 356 15210 412 15219
rect 0 15113 28 15161
rect 356 15038 412 15047
rect 356 14973 412 14982
rect 0 14859 28 14907
rect 356 14801 412 14810
rect 356 14736 412 14745
rect 0 14639 28 14687
rect 0 14543 28 14591
rect 356 14485 412 14494
rect 356 14420 412 14429
rect 0 14323 28 14371
rect 356 14248 412 14257
rect 356 14183 412 14192
rect 0 14069 28 14117
rect 356 14011 412 14020
rect 356 13946 412 13955
rect 0 13849 28 13897
rect 0 13753 28 13801
rect 356 13695 412 13704
rect 356 13630 412 13639
rect 0 13533 28 13581
rect 356 13458 412 13467
rect 356 13393 412 13402
rect 0 13279 28 13327
rect 356 13221 412 13230
rect 356 13156 412 13165
rect 0 13059 28 13107
rect 0 12963 28 13011
rect 356 12905 412 12914
rect 356 12840 412 12849
rect 0 12743 28 12791
rect 356 12668 412 12677
rect 356 12603 412 12612
rect 0 12489 28 12537
rect 356 12431 412 12440
rect 356 12366 412 12375
rect 0 12269 28 12317
rect 0 12173 28 12221
rect 356 12115 412 12124
rect 356 12050 412 12059
rect 0 11953 28 12001
rect 356 11878 412 11887
rect 356 11813 412 11822
rect 0 11699 28 11747
rect 356 11641 412 11650
rect 356 11576 412 11585
rect 0 11479 28 11527
rect 0 11383 28 11431
rect 356 11325 412 11334
rect 356 11260 412 11269
rect 0 11163 28 11211
rect 356 11088 412 11097
rect 356 11023 412 11032
rect 0 10909 28 10957
rect 356 10851 412 10860
rect 356 10786 412 10795
rect 0 10689 28 10737
rect 0 10593 28 10641
rect 356 10535 412 10544
rect 356 10470 412 10479
rect 0 10373 28 10421
rect 356 10298 412 10307
rect 356 10233 412 10242
rect 0 10119 28 10167
rect 356 10061 412 10070
rect 356 9996 412 10005
rect 0 9899 28 9947
rect 0 9803 28 9851
rect 356 9745 412 9754
rect 356 9680 412 9689
rect 0 9583 28 9631
rect 356 9508 412 9517
rect 356 9443 412 9452
rect 0 9329 28 9377
rect 356 9271 412 9280
rect 356 9206 412 9215
rect 0 9109 28 9157
rect 0 9013 28 9061
rect 356 8955 412 8964
rect 356 8890 412 8899
rect 0 8793 28 8841
rect 356 8718 412 8727
rect 356 8653 412 8662
rect 0 8539 28 8587
rect 356 8481 412 8490
rect 356 8416 412 8425
rect 0 8319 28 8367
rect 0 8223 28 8271
rect 356 8165 412 8174
rect 356 8100 412 8109
rect 0 8003 28 8051
rect 356 7928 412 7937
rect 356 7863 412 7872
rect 0 7749 28 7797
rect 356 7691 412 7700
rect 356 7626 412 7635
rect 0 7529 28 7577
rect 0 7433 28 7481
rect 356 7375 412 7384
rect 356 7310 412 7319
rect 0 7213 28 7261
rect 356 7138 412 7147
rect 356 7073 412 7082
rect 0 6959 28 7007
rect 356 6901 412 6910
rect 356 6836 412 6845
rect 0 6739 28 6787
rect 0 6643 28 6691
rect 356 6585 412 6594
rect 356 6520 412 6529
rect 0 6423 28 6471
rect 356 6348 412 6357
rect 356 6283 412 6292
rect 0 6169 28 6217
rect 356 6111 412 6120
rect 356 6046 412 6055
rect 0 5949 28 5997
rect 0 5853 28 5901
rect 356 5795 412 5804
rect 356 5730 412 5739
rect 0 5633 28 5681
rect 356 5558 412 5567
rect 356 5493 412 5502
rect 0 5379 28 5427
rect 356 5321 412 5330
rect 356 5256 412 5265
rect 0 5159 28 5207
rect 0 5063 28 5111
rect 356 5005 412 5014
rect 356 4940 412 4949
rect 0 4843 28 4891
rect 356 4768 412 4777
rect 356 4703 412 4712
rect 0 4589 28 4637
rect 356 4531 412 4540
rect 356 4466 412 4475
rect 0 4369 28 4417
rect 0 4273 28 4321
rect 356 4215 412 4224
rect 356 4150 412 4159
rect 0 4053 28 4101
rect 356 3978 412 3987
rect 356 3913 412 3922
rect 0 3799 28 3847
rect 356 3741 412 3750
rect 356 3676 412 3685
rect 0 3579 28 3627
rect 0 3483 28 3531
rect 356 3425 412 3434
rect 356 3360 412 3369
rect 0 3263 28 3311
rect 356 3188 412 3197
rect 356 3123 412 3132
rect 0 3009 28 3057
rect 356 2951 412 2960
rect 356 2886 412 2895
rect 0 2789 28 2837
rect 0 2693 28 2741
rect 356 2635 412 2644
rect 356 2570 412 2579
rect 0 2473 28 2521
rect 356 2398 412 2407
rect 356 2333 412 2342
rect 0 2219 28 2267
rect 356 2161 412 2170
rect 356 2096 412 2105
rect 0 1999 28 2047
rect 0 1903 28 1951
rect 356 1845 412 1854
rect 356 1780 412 1789
rect 0 1683 28 1731
rect 356 1608 412 1617
rect 356 1543 412 1552
rect 0 1429 28 1477
rect 356 1371 412 1380
rect 356 1306 412 1315
rect 0 1209 28 1257
rect 0 1113 28 1161
rect 356 1055 412 1064
rect 356 990 412 999
rect 0 893 28 941
rect 356 818 412 827
rect 356 753 412 762
<< via2 >>
rect 356 51322 412 51378
rect 356 51085 412 51141
rect 356 50769 412 50825
rect 356 50532 412 50588
rect 356 50295 412 50351
rect 356 49979 412 50035
rect 356 49742 412 49798
rect 356 49505 412 49561
rect 356 49189 412 49245
rect 356 48952 412 49008
rect 356 48715 412 48771
rect 356 48399 412 48455
rect 356 48162 412 48218
rect 356 47925 412 47981
rect 356 47609 412 47665
rect 356 47372 412 47428
rect 356 47135 412 47191
rect 356 46819 412 46875
rect 356 46582 412 46638
rect 356 46345 412 46401
rect 356 46029 412 46085
rect 356 45792 412 45848
rect 356 45555 412 45611
rect 356 45239 412 45295
rect 356 45002 412 45058
rect 356 44765 412 44821
rect 356 44449 412 44505
rect 356 44212 412 44268
rect 356 43975 412 44031
rect 356 43659 412 43715
rect 356 43422 412 43478
rect 356 43185 412 43241
rect 356 42869 412 42925
rect 356 42632 412 42688
rect 356 42395 412 42451
rect 356 42079 412 42135
rect 356 41842 412 41898
rect 356 41605 412 41661
rect 356 41289 412 41345
rect 356 41052 412 41108
rect 356 40815 412 40871
rect 356 40499 412 40555
rect 356 40262 412 40318
rect 356 40025 412 40081
rect 356 39709 412 39765
rect 356 39472 412 39528
rect 356 39235 412 39291
rect 356 38919 412 38975
rect 356 38682 412 38738
rect 356 38445 412 38501
rect 356 38129 412 38185
rect 356 37892 412 37948
rect 356 37655 412 37711
rect 356 37339 412 37395
rect 356 37102 412 37158
rect 356 36865 412 36921
rect 356 36549 412 36605
rect 356 36312 412 36368
rect 356 36075 412 36131
rect 356 35759 412 35815
rect 356 35522 412 35578
rect 356 35285 412 35341
rect 356 34969 412 35025
rect 356 34732 412 34788
rect 356 34495 412 34551
rect 356 34179 412 34235
rect 356 33942 412 33998
rect 356 33705 412 33761
rect 356 33389 412 33445
rect 356 33152 412 33208
rect 356 32915 412 32971
rect 356 32599 412 32655
rect 356 32362 412 32418
rect 356 32125 412 32181
rect 356 31809 412 31865
rect 356 31572 412 31628
rect 356 31335 412 31391
rect 356 31019 412 31075
rect 356 30782 412 30838
rect 356 30545 412 30601
rect 356 30229 412 30285
rect 356 29992 412 30048
rect 356 29755 412 29811
rect 356 29439 412 29495
rect 356 29202 412 29258
rect 356 28965 412 29021
rect 356 28649 412 28705
rect 356 28412 412 28468
rect 356 28175 412 28231
rect 356 27859 412 27915
rect 356 27622 412 27678
rect 356 27385 412 27441
rect 356 27069 412 27125
rect 356 26832 412 26888
rect 356 26595 412 26651
rect 356 26279 412 26335
rect 356 26042 412 26098
rect 356 25805 412 25861
rect 356 25489 412 25545
rect 356 25252 412 25308
rect 356 25015 412 25071
rect 356 24699 412 24755
rect 356 24462 412 24518
rect 356 24225 412 24281
rect 356 23909 412 23965
rect 356 23672 412 23728
rect 356 23435 412 23491
rect 356 23119 412 23175
rect 356 22882 412 22938
rect 356 22645 412 22701
rect 356 22329 412 22385
rect 356 22092 412 22148
rect 356 21855 412 21911
rect 356 21539 412 21595
rect 356 21302 412 21358
rect 356 21065 412 21121
rect 356 20749 412 20805
rect 356 20512 412 20568
rect 356 20275 412 20331
rect 356 19959 412 20015
rect 356 19722 412 19778
rect 356 19485 412 19541
rect 356 19169 412 19225
rect 356 18932 412 18988
rect 356 18695 412 18751
rect 356 18379 412 18435
rect 356 18142 412 18198
rect 356 17905 412 17961
rect 356 17589 412 17645
rect 356 17352 412 17408
rect 356 17115 412 17171
rect 356 16799 412 16855
rect 356 16562 412 16618
rect 356 16325 412 16381
rect 356 16009 412 16065
rect 356 15772 412 15828
rect 356 15535 412 15591
rect 356 15219 412 15275
rect 356 14982 412 15038
rect 356 14745 412 14801
rect 356 14429 412 14485
rect 356 14192 412 14248
rect 356 13955 412 14011
rect 356 13639 412 13695
rect 356 13402 412 13458
rect 356 13165 412 13221
rect 356 12849 412 12905
rect 356 12612 412 12668
rect 356 12375 412 12431
rect 356 12059 412 12115
rect 356 11822 412 11878
rect 356 11585 412 11641
rect 356 11269 412 11325
rect 356 11032 412 11088
rect 356 10795 412 10851
rect 356 10479 412 10535
rect 356 10242 412 10298
rect 356 10005 412 10061
rect 356 9689 412 9745
rect 356 9452 412 9508
rect 356 9215 412 9271
rect 356 8899 412 8955
rect 356 8662 412 8718
rect 356 8425 412 8481
rect 356 8109 412 8165
rect 356 7872 412 7928
rect 356 7635 412 7691
rect 356 7319 412 7375
rect 356 7082 412 7138
rect 356 6845 412 6901
rect 356 6529 412 6585
rect 356 6292 412 6348
rect 356 6055 412 6111
rect 356 5739 412 5795
rect 356 5502 412 5558
rect 356 5265 412 5321
rect 356 4949 412 5005
rect 356 4712 412 4768
rect 356 4475 412 4531
rect 356 4159 412 4215
rect 356 3922 412 3978
rect 356 3685 412 3741
rect 356 3369 412 3425
rect 356 3132 412 3188
rect 356 2895 412 2951
rect 356 2579 412 2635
rect 356 2342 412 2398
rect 356 2105 412 2161
rect 356 1789 412 1845
rect 356 1552 412 1608
rect 356 1315 412 1371
rect 356 999 412 1055
rect 356 762 412 818
<< metal3 >>
rect 335 51378 433 51399
rect 335 51322 356 51378
rect 412 51322 433 51378
rect 335 51301 433 51322
rect 335 51141 433 51162
rect 335 51085 356 51141
rect 412 51085 433 51141
rect 335 51064 433 51085
rect 335 50825 433 50846
rect 335 50769 356 50825
rect 412 50769 433 50825
rect 335 50748 433 50769
rect 335 50588 433 50609
rect 335 50532 356 50588
rect 412 50532 433 50588
rect 335 50511 433 50532
rect 335 50351 433 50372
rect 335 50295 356 50351
rect 412 50295 433 50351
rect 335 50274 433 50295
rect 335 50035 433 50056
rect 335 49979 356 50035
rect 412 49979 433 50035
rect 335 49958 433 49979
rect 335 49798 433 49819
rect 335 49742 356 49798
rect 412 49742 433 49798
rect 335 49721 433 49742
rect 335 49561 433 49582
rect 335 49505 356 49561
rect 412 49505 433 49561
rect 335 49484 433 49505
rect 335 49245 433 49266
rect 335 49189 356 49245
rect 412 49189 433 49245
rect 335 49168 433 49189
rect 335 49008 433 49029
rect 335 48952 356 49008
rect 412 48952 433 49008
rect 335 48931 433 48952
rect 335 48771 433 48792
rect 335 48715 356 48771
rect 412 48715 433 48771
rect 335 48694 433 48715
rect 335 48455 433 48476
rect 335 48399 356 48455
rect 412 48399 433 48455
rect 335 48378 433 48399
rect 335 48218 433 48239
rect 335 48162 356 48218
rect 412 48162 433 48218
rect 335 48141 433 48162
rect 335 47981 433 48002
rect 335 47925 356 47981
rect 412 47925 433 47981
rect 335 47904 433 47925
rect 335 47665 433 47686
rect 335 47609 356 47665
rect 412 47609 433 47665
rect 335 47588 433 47609
rect 335 47428 433 47449
rect 335 47372 356 47428
rect 412 47372 433 47428
rect 335 47351 433 47372
rect 335 47191 433 47212
rect 335 47135 356 47191
rect 412 47135 433 47191
rect 335 47114 433 47135
rect 335 46875 433 46896
rect 335 46819 356 46875
rect 412 46819 433 46875
rect 335 46798 433 46819
rect 335 46638 433 46659
rect 335 46582 356 46638
rect 412 46582 433 46638
rect 335 46561 433 46582
rect 335 46401 433 46422
rect 335 46345 356 46401
rect 412 46345 433 46401
rect 335 46324 433 46345
rect 335 46085 433 46106
rect 335 46029 356 46085
rect 412 46029 433 46085
rect 335 46008 433 46029
rect 335 45848 433 45869
rect 335 45792 356 45848
rect 412 45792 433 45848
rect 335 45771 433 45792
rect 335 45611 433 45632
rect 335 45555 356 45611
rect 412 45555 433 45611
rect 335 45534 433 45555
rect 335 45295 433 45316
rect 335 45239 356 45295
rect 412 45239 433 45295
rect 335 45218 433 45239
rect 335 45058 433 45079
rect 335 45002 356 45058
rect 412 45002 433 45058
rect 335 44981 433 45002
rect 335 44821 433 44842
rect 335 44765 356 44821
rect 412 44765 433 44821
rect 335 44744 433 44765
rect 335 44505 433 44526
rect 335 44449 356 44505
rect 412 44449 433 44505
rect 335 44428 433 44449
rect 335 44268 433 44289
rect 335 44212 356 44268
rect 412 44212 433 44268
rect 335 44191 433 44212
rect 335 44031 433 44052
rect 335 43975 356 44031
rect 412 43975 433 44031
rect 335 43954 433 43975
rect 335 43715 433 43736
rect 335 43659 356 43715
rect 412 43659 433 43715
rect 335 43638 433 43659
rect 335 43478 433 43499
rect 335 43422 356 43478
rect 412 43422 433 43478
rect 335 43401 433 43422
rect 335 43241 433 43262
rect 335 43185 356 43241
rect 412 43185 433 43241
rect 335 43164 433 43185
rect 335 42925 433 42946
rect 335 42869 356 42925
rect 412 42869 433 42925
rect 335 42848 433 42869
rect 335 42688 433 42709
rect 335 42632 356 42688
rect 412 42632 433 42688
rect 335 42611 433 42632
rect 335 42451 433 42472
rect 335 42395 356 42451
rect 412 42395 433 42451
rect 335 42374 433 42395
rect 335 42135 433 42156
rect 335 42079 356 42135
rect 412 42079 433 42135
rect 335 42058 433 42079
rect 335 41898 433 41919
rect 335 41842 356 41898
rect 412 41842 433 41898
rect 335 41821 433 41842
rect 335 41661 433 41682
rect 335 41605 356 41661
rect 412 41605 433 41661
rect 335 41584 433 41605
rect 335 41345 433 41366
rect 335 41289 356 41345
rect 412 41289 433 41345
rect 335 41268 433 41289
rect 335 41108 433 41129
rect 335 41052 356 41108
rect 412 41052 433 41108
rect 335 41031 433 41052
rect 335 40871 433 40892
rect 335 40815 356 40871
rect 412 40815 433 40871
rect 335 40794 433 40815
rect 335 40555 433 40576
rect 335 40499 356 40555
rect 412 40499 433 40555
rect 335 40478 433 40499
rect 335 40318 433 40339
rect 335 40262 356 40318
rect 412 40262 433 40318
rect 335 40241 433 40262
rect 335 40081 433 40102
rect 335 40025 356 40081
rect 412 40025 433 40081
rect 335 40004 433 40025
rect 335 39765 433 39786
rect 335 39709 356 39765
rect 412 39709 433 39765
rect 335 39688 433 39709
rect 335 39528 433 39549
rect 335 39472 356 39528
rect 412 39472 433 39528
rect 335 39451 433 39472
rect 335 39291 433 39312
rect 335 39235 356 39291
rect 412 39235 433 39291
rect 335 39214 433 39235
rect 335 38975 433 38996
rect 335 38919 356 38975
rect 412 38919 433 38975
rect 335 38898 433 38919
rect 335 38738 433 38759
rect 335 38682 356 38738
rect 412 38682 433 38738
rect 335 38661 433 38682
rect 335 38501 433 38522
rect 335 38445 356 38501
rect 412 38445 433 38501
rect 335 38424 433 38445
rect 335 38185 433 38206
rect 335 38129 356 38185
rect 412 38129 433 38185
rect 335 38108 433 38129
rect 335 37948 433 37969
rect 335 37892 356 37948
rect 412 37892 433 37948
rect 335 37871 433 37892
rect 335 37711 433 37732
rect 335 37655 356 37711
rect 412 37655 433 37711
rect 335 37634 433 37655
rect 335 37395 433 37416
rect 335 37339 356 37395
rect 412 37339 433 37395
rect 335 37318 433 37339
rect 335 37158 433 37179
rect 335 37102 356 37158
rect 412 37102 433 37158
rect 335 37081 433 37102
rect 335 36921 433 36942
rect 335 36865 356 36921
rect 412 36865 433 36921
rect 335 36844 433 36865
rect 335 36605 433 36626
rect 335 36549 356 36605
rect 412 36549 433 36605
rect 335 36528 433 36549
rect 335 36368 433 36389
rect 335 36312 356 36368
rect 412 36312 433 36368
rect 335 36291 433 36312
rect 335 36131 433 36152
rect 335 36075 356 36131
rect 412 36075 433 36131
rect 335 36054 433 36075
rect 335 35815 433 35836
rect 335 35759 356 35815
rect 412 35759 433 35815
rect 335 35738 433 35759
rect 335 35578 433 35599
rect 335 35522 356 35578
rect 412 35522 433 35578
rect 335 35501 433 35522
rect 335 35341 433 35362
rect 335 35285 356 35341
rect 412 35285 433 35341
rect 335 35264 433 35285
rect 335 35025 433 35046
rect 335 34969 356 35025
rect 412 34969 433 35025
rect 335 34948 433 34969
rect 335 34788 433 34809
rect 335 34732 356 34788
rect 412 34732 433 34788
rect 335 34711 433 34732
rect 335 34551 433 34572
rect 335 34495 356 34551
rect 412 34495 433 34551
rect 335 34474 433 34495
rect 335 34235 433 34256
rect 335 34179 356 34235
rect 412 34179 433 34235
rect 335 34158 433 34179
rect 335 33998 433 34019
rect 335 33942 356 33998
rect 412 33942 433 33998
rect 335 33921 433 33942
rect 335 33761 433 33782
rect 335 33705 356 33761
rect 412 33705 433 33761
rect 335 33684 433 33705
rect 335 33445 433 33466
rect 335 33389 356 33445
rect 412 33389 433 33445
rect 335 33368 433 33389
rect 335 33208 433 33229
rect 335 33152 356 33208
rect 412 33152 433 33208
rect 335 33131 433 33152
rect 335 32971 433 32992
rect 335 32915 356 32971
rect 412 32915 433 32971
rect 335 32894 433 32915
rect 335 32655 433 32676
rect 335 32599 356 32655
rect 412 32599 433 32655
rect 335 32578 433 32599
rect 335 32418 433 32439
rect 335 32362 356 32418
rect 412 32362 433 32418
rect 335 32341 433 32362
rect 335 32181 433 32202
rect 335 32125 356 32181
rect 412 32125 433 32181
rect 335 32104 433 32125
rect 335 31865 433 31886
rect 335 31809 356 31865
rect 412 31809 433 31865
rect 335 31788 433 31809
rect 335 31628 433 31649
rect 335 31572 356 31628
rect 412 31572 433 31628
rect 335 31551 433 31572
rect 335 31391 433 31412
rect 335 31335 356 31391
rect 412 31335 433 31391
rect 335 31314 433 31335
rect 335 31075 433 31096
rect 335 31019 356 31075
rect 412 31019 433 31075
rect 335 30998 433 31019
rect 335 30838 433 30859
rect 335 30782 356 30838
rect 412 30782 433 30838
rect 335 30761 433 30782
rect 335 30601 433 30622
rect 335 30545 356 30601
rect 412 30545 433 30601
rect 335 30524 433 30545
rect 335 30285 433 30306
rect 335 30229 356 30285
rect 412 30229 433 30285
rect 335 30208 433 30229
rect 335 30048 433 30069
rect 335 29992 356 30048
rect 412 29992 433 30048
rect 335 29971 433 29992
rect 335 29811 433 29832
rect 335 29755 356 29811
rect 412 29755 433 29811
rect 335 29734 433 29755
rect 335 29495 433 29516
rect 335 29439 356 29495
rect 412 29439 433 29495
rect 335 29418 433 29439
rect 335 29258 433 29279
rect 335 29202 356 29258
rect 412 29202 433 29258
rect 335 29181 433 29202
rect 335 29021 433 29042
rect 335 28965 356 29021
rect 412 28965 433 29021
rect 335 28944 433 28965
rect 335 28705 433 28726
rect 335 28649 356 28705
rect 412 28649 433 28705
rect 335 28628 433 28649
rect 335 28468 433 28489
rect 335 28412 356 28468
rect 412 28412 433 28468
rect 335 28391 433 28412
rect 335 28231 433 28252
rect 335 28175 356 28231
rect 412 28175 433 28231
rect 335 28154 433 28175
rect 335 27915 433 27936
rect 335 27859 356 27915
rect 412 27859 433 27915
rect 335 27838 433 27859
rect 335 27678 433 27699
rect 335 27622 356 27678
rect 412 27622 433 27678
rect 335 27601 433 27622
rect 335 27441 433 27462
rect 335 27385 356 27441
rect 412 27385 433 27441
rect 335 27364 433 27385
rect 335 27125 433 27146
rect 335 27069 356 27125
rect 412 27069 433 27125
rect 335 27048 433 27069
rect 335 26888 433 26909
rect 335 26832 356 26888
rect 412 26832 433 26888
rect 335 26811 433 26832
rect 335 26651 433 26672
rect 335 26595 356 26651
rect 412 26595 433 26651
rect 335 26574 433 26595
rect 335 26335 433 26356
rect 335 26279 356 26335
rect 412 26279 433 26335
rect 335 26258 433 26279
rect 335 26098 433 26119
rect 335 26042 356 26098
rect 412 26042 433 26098
rect 335 26021 433 26042
rect 335 25861 433 25882
rect 335 25805 356 25861
rect 412 25805 433 25861
rect 335 25784 433 25805
rect 335 25545 433 25566
rect 335 25489 356 25545
rect 412 25489 433 25545
rect 335 25468 433 25489
rect 335 25308 433 25329
rect 335 25252 356 25308
rect 412 25252 433 25308
rect 335 25231 433 25252
rect 335 25071 433 25092
rect 335 25015 356 25071
rect 412 25015 433 25071
rect 335 24994 433 25015
rect 335 24755 433 24776
rect 335 24699 356 24755
rect 412 24699 433 24755
rect 335 24678 433 24699
rect 335 24518 433 24539
rect 335 24462 356 24518
rect 412 24462 433 24518
rect 335 24441 433 24462
rect 335 24281 433 24302
rect 335 24225 356 24281
rect 412 24225 433 24281
rect 335 24204 433 24225
rect 335 23965 433 23986
rect 335 23909 356 23965
rect 412 23909 433 23965
rect 335 23888 433 23909
rect 335 23728 433 23749
rect 335 23672 356 23728
rect 412 23672 433 23728
rect 335 23651 433 23672
rect 335 23491 433 23512
rect 335 23435 356 23491
rect 412 23435 433 23491
rect 335 23414 433 23435
rect 335 23175 433 23196
rect 335 23119 356 23175
rect 412 23119 433 23175
rect 335 23098 433 23119
rect 335 22938 433 22959
rect 335 22882 356 22938
rect 412 22882 433 22938
rect 335 22861 433 22882
rect 335 22701 433 22722
rect 335 22645 356 22701
rect 412 22645 433 22701
rect 335 22624 433 22645
rect 335 22385 433 22406
rect 335 22329 356 22385
rect 412 22329 433 22385
rect 335 22308 433 22329
rect 335 22148 433 22169
rect 335 22092 356 22148
rect 412 22092 433 22148
rect 335 22071 433 22092
rect 335 21911 433 21932
rect 335 21855 356 21911
rect 412 21855 433 21911
rect 335 21834 433 21855
rect 335 21595 433 21616
rect 335 21539 356 21595
rect 412 21539 433 21595
rect 335 21518 433 21539
rect 335 21358 433 21379
rect 335 21302 356 21358
rect 412 21302 433 21358
rect 335 21281 433 21302
rect 335 21121 433 21142
rect 335 21065 356 21121
rect 412 21065 433 21121
rect 335 21044 433 21065
rect 335 20805 433 20826
rect 335 20749 356 20805
rect 412 20749 433 20805
rect 335 20728 433 20749
rect 335 20568 433 20589
rect 335 20512 356 20568
rect 412 20512 433 20568
rect 335 20491 433 20512
rect 335 20331 433 20352
rect 335 20275 356 20331
rect 412 20275 433 20331
rect 335 20254 433 20275
rect 335 20015 433 20036
rect 335 19959 356 20015
rect 412 19959 433 20015
rect 335 19938 433 19959
rect 335 19778 433 19799
rect 335 19722 356 19778
rect 412 19722 433 19778
rect 335 19701 433 19722
rect 335 19541 433 19562
rect 335 19485 356 19541
rect 412 19485 433 19541
rect 335 19464 433 19485
rect 335 19225 433 19246
rect 335 19169 356 19225
rect 412 19169 433 19225
rect 335 19148 433 19169
rect 335 18988 433 19009
rect 335 18932 356 18988
rect 412 18932 433 18988
rect 335 18911 433 18932
rect 335 18751 433 18772
rect 335 18695 356 18751
rect 412 18695 433 18751
rect 335 18674 433 18695
rect 335 18435 433 18456
rect 335 18379 356 18435
rect 412 18379 433 18435
rect 335 18358 433 18379
rect 335 18198 433 18219
rect 335 18142 356 18198
rect 412 18142 433 18198
rect 335 18121 433 18142
rect 335 17961 433 17982
rect 335 17905 356 17961
rect 412 17905 433 17961
rect 335 17884 433 17905
rect 335 17645 433 17666
rect 335 17589 356 17645
rect 412 17589 433 17645
rect 335 17568 433 17589
rect 335 17408 433 17429
rect 335 17352 356 17408
rect 412 17352 433 17408
rect 335 17331 433 17352
rect 335 17171 433 17192
rect 335 17115 356 17171
rect 412 17115 433 17171
rect 335 17094 433 17115
rect 335 16855 433 16876
rect 335 16799 356 16855
rect 412 16799 433 16855
rect 335 16778 433 16799
rect 335 16618 433 16639
rect 335 16562 356 16618
rect 412 16562 433 16618
rect 335 16541 433 16562
rect 335 16381 433 16402
rect 335 16325 356 16381
rect 412 16325 433 16381
rect 335 16304 433 16325
rect 335 16065 433 16086
rect 335 16009 356 16065
rect 412 16009 433 16065
rect 335 15988 433 16009
rect 335 15828 433 15849
rect 335 15772 356 15828
rect 412 15772 433 15828
rect 335 15751 433 15772
rect 335 15591 433 15612
rect 335 15535 356 15591
rect 412 15535 433 15591
rect 335 15514 433 15535
rect 335 15275 433 15296
rect 335 15219 356 15275
rect 412 15219 433 15275
rect 335 15198 433 15219
rect 335 15038 433 15059
rect 335 14982 356 15038
rect 412 14982 433 15038
rect 335 14961 433 14982
rect 335 14801 433 14822
rect 335 14745 356 14801
rect 412 14745 433 14801
rect 335 14724 433 14745
rect 335 14485 433 14506
rect 335 14429 356 14485
rect 412 14429 433 14485
rect 335 14408 433 14429
rect 335 14248 433 14269
rect 335 14192 356 14248
rect 412 14192 433 14248
rect 335 14171 433 14192
rect 335 14011 433 14032
rect 335 13955 356 14011
rect 412 13955 433 14011
rect 335 13934 433 13955
rect 335 13695 433 13716
rect 335 13639 356 13695
rect 412 13639 433 13695
rect 335 13618 433 13639
rect 335 13458 433 13479
rect 335 13402 356 13458
rect 412 13402 433 13458
rect 335 13381 433 13402
rect 335 13221 433 13242
rect 335 13165 356 13221
rect 412 13165 433 13221
rect 335 13144 433 13165
rect 335 12905 433 12926
rect 335 12849 356 12905
rect 412 12849 433 12905
rect 335 12828 433 12849
rect 335 12668 433 12689
rect 335 12612 356 12668
rect 412 12612 433 12668
rect 335 12591 433 12612
rect 335 12431 433 12452
rect 335 12375 356 12431
rect 412 12375 433 12431
rect 335 12354 433 12375
rect 335 12115 433 12136
rect 335 12059 356 12115
rect 412 12059 433 12115
rect 335 12038 433 12059
rect 335 11878 433 11899
rect 335 11822 356 11878
rect 412 11822 433 11878
rect 335 11801 433 11822
rect 335 11641 433 11662
rect 335 11585 356 11641
rect 412 11585 433 11641
rect 335 11564 433 11585
rect 335 11325 433 11346
rect 335 11269 356 11325
rect 412 11269 433 11325
rect 335 11248 433 11269
rect 335 11088 433 11109
rect 335 11032 356 11088
rect 412 11032 433 11088
rect 335 11011 433 11032
rect 335 10851 433 10872
rect 335 10795 356 10851
rect 412 10795 433 10851
rect 335 10774 433 10795
rect 335 10535 433 10556
rect 335 10479 356 10535
rect 412 10479 433 10535
rect 335 10458 433 10479
rect 335 10298 433 10319
rect 335 10242 356 10298
rect 412 10242 433 10298
rect 335 10221 433 10242
rect 335 10061 433 10082
rect 335 10005 356 10061
rect 412 10005 433 10061
rect 335 9984 433 10005
rect 335 9745 433 9766
rect 335 9689 356 9745
rect 412 9689 433 9745
rect 335 9668 433 9689
rect 335 9508 433 9529
rect 335 9452 356 9508
rect 412 9452 433 9508
rect 335 9431 433 9452
rect 335 9271 433 9292
rect 335 9215 356 9271
rect 412 9215 433 9271
rect 335 9194 433 9215
rect 335 8955 433 8976
rect 335 8899 356 8955
rect 412 8899 433 8955
rect 335 8878 433 8899
rect 335 8718 433 8739
rect 335 8662 356 8718
rect 412 8662 433 8718
rect 335 8641 433 8662
rect 335 8481 433 8502
rect 335 8425 356 8481
rect 412 8425 433 8481
rect 335 8404 433 8425
rect 335 8165 433 8186
rect 335 8109 356 8165
rect 412 8109 433 8165
rect 335 8088 433 8109
rect 335 7928 433 7949
rect 335 7872 356 7928
rect 412 7872 433 7928
rect 335 7851 433 7872
rect 335 7691 433 7712
rect 335 7635 356 7691
rect 412 7635 433 7691
rect 335 7614 433 7635
rect 335 7375 433 7396
rect 335 7319 356 7375
rect 412 7319 433 7375
rect 335 7298 433 7319
rect 335 7138 433 7159
rect 335 7082 356 7138
rect 412 7082 433 7138
rect 335 7061 433 7082
rect 335 6901 433 6922
rect 335 6845 356 6901
rect 412 6845 433 6901
rect 335 6824 433 6845
rect 335 6585 433 6606
rect 335 6529 356 6585
rect 412 6529 433 6585
rect 335 6508 433 6529
rect 335 6348 433 6369
rect 335 6292 356 6348
rect 412 6292 433 6348
rect 335 6271 433 6292
rect 335 6111 433 6132
rect 335 6055 356 6111
rect 412 6055 433 6111
rect 335 6034 433 6055
rect 335 5795 433 5816
rect 335 5739 356 5795
rect 412 5739 433 5795
rect 335 5718 433 5739
rect 335 5558 433 5579
rect 335 5502 356 5558
rect 412 5502 433 5558
rect 335 5481 433 5502
rect 335 5321 433 5342
rect 335 5265 356 5321
rect 412 5265 433 5321
rect 335 5244 433 5265
rect 335 5005 433 5026
rect 335 4949 356 5005
rect 412 4949 433 5005
rect 335 4928 433 4949
rect 335 4768 433 4789
rect 335 4712 356 4768
rect 412 4712 433 4768
rect 335 4691 433 4712
rect 335 4531 433 4552
rect 335 4475 356 4531
rect 412 4475 433 4531
rect 335 4454 433 4475
rect 335 4215 433 4236
rect 335 4159 356 4215
rect 412 4159 433 4215
rect 335 4138 433 4159
rect 335 3978 433 3999
rect 335 3922 356 3978
rect 412 3922 433 3978
rect 335 3901 433 3922
rect 335 3741 433 3762
rect 335 3685 356 3741
rect 412 3685 433 3741
rect 335 3664 433 3685
rect 335 3425 433 3446
rect 335 3369 356 3425
rect 412 3369 433 3425
rect 335 3348 433 3369
rect 335 3188 433 3209
rect 335 3132 356 3188
rect 412 3132 433 3188
rect 335 3111 433 3132
rect 335 2951 433 2972
rect 335 2895 356 2951
rect 412 2895 433 2951
rect 335 2874 433 2895
rect 335 2635 433 2656
rect 335 2579 356 2635
rect 412 2579 433 2635
rect 335 2558 433 2579
rect 335 2398 433 2419
rect 335 2342 356 2398
rect 412 2342 433 2398
rect 335 2321 433 2342
rect 335 2161 433 2182
rect 335 2105 356 2161
rect 412 2105 433 2161
rect 335 2084 433 2105
rect 335 1845 433 1866
rect 335 1789 356 1845
rect 412 1789 433 1845
rect 335 1768 433 1789
rect 335 1608 433 1629
rect 335 1552 356 1608
rect 412 1552 433 1608
rect 335 1531 433 1552
rect 335 1371 433 1392
rect 335 1315 356 1371
rect 412 1315 433 1371
rect 335 1294 433 1315
rect 335 1055 433 1076
rect 335 999 356 1055
rect 412 999 433 1055
rect 335 978 433 999
rect 335 818 433 839
rect 335 762 356 818
rect 412 762 433 818
rect 335 741 433 762
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_0
timestamp 1723858470
transform -1 0 624 0 -1 3160
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_1
timestamp 1723858470
transform -1 0 624 0 1 2370
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_2
timestamp 1723858470
transform -1 0 624 0 -1 2370
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_3
timestamp 1723858470
transform -1 0 624 0 1 790
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_4
timestamp 1723858470
transform -1 0 624 0 -1 790
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_5
timestamp 1723858470
transform -1 0 624 0 1 1580
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_6
timestamp 1723858470
transform -1 0 624 0 -1 1580
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_7
timestamp 1723858470
transform -1 0 624 0 1 12640
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_8
timestamp 1723858470
transform -1 0 624 0 -1 12640
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_9
timestamp 1723858470
transform -1 0 624 0 1 11850
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_10
timestamp 1723858470
transform -1 0 624 0 -1 11850
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_11
timestamp 1723858470
transform -1 0 624 0 1 11060
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_12
timestamp 1723858470
transform -1 0 624 0 -1 11060
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_13
timestamp 1723858470
transform -1 0 624 0 1 10270
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_14
timestamp 1723858470
transform -1 0 624 0 -1 10270
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_15
timestamp 1723858470
transform -1 0 624 0 1 9480
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_16
timestamp 1723858470
transform -1 0 624 0 -1 9480
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_17
timestamp 1723858470
transform -1 0 624 0 1 8690
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_18
timestamp 1723858470
transform -1 0 624 0 -1 8690
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_19
timestamp 1723858470
transform -1 0 624 0 1 7900
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_20
timestamp 1723858470
transform -1 0 624 0 -1 7900
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_21
timestamp 1723858470
transform -1 0 624 0 1 7110
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_22
timestamp 1723858470
transform -1 0 624 0 -1 7110
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_23
timestamp 1723858470
transform -1 0 624 0 1 6320
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_24
timestamp 1723858470
transform -1 0 624 0 -1 6320
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_25
timestamp 1723858470
transform -1 0 624 0 1 5530
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_26
timestamp 1723858470
transform -1 0 624 0 -1 5530
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_27
timestamp 1723858470
transform -1 0 624 0 1 4740
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_28
timestamp 1723858470
transform -1 0 624 0 -1 4740
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_29
timestamp 1723858470
transform -1 0 624 0 1 3950
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_30
timestamp 1723858470
transform -1 0 624 0 -1 3950
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_31
timestamp 1723858470
transform -1 0 624 0 1 3160
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_32
timestamp 1723858470
transform -1 0 624 0 1 25280
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_33
timestamp 1723858470
transform -1 0 624 0 -1 25280
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_34
timestamp 1723858470
transform -1 0 624 0 1 24490
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_35
timestamp 1723858470
transform -1 0 624 0 -1 24490
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_36
timestamp 1723858470
transform -1 0 624 0 1 23700
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_37
timestamp 1723858470
transform -1 0 624 0 -1 23700
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_38
timestamp 1723858470
transform -1 0 624 0 1 22910
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_39
timestamp 1723858470
transform -1 0 624 0 -1 22910
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_40
timestamp 1723858470
transform -1 0 624 0 1 22120
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_41
timestamp 1723858470
transform -1 0 624 0 -1 22120
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_42
timestamp 1723858470
transform -1 0 624 0 1 21330
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_43
timestamp 1723858470
transform -1 0 624 0 -1 21330
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_44
timestamp 1723858470
transform -1 0 624 0 1 20540
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_45
timestamp 1723858470
transform -1 0 624 0 -1 20540
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_46
timestamp 1723858470
transform -1 0 624 0 1 19750
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_47
timestamp 1723858470
transform -1 0 624 0 -1 19750
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_48
timestamp 1723858470
transform -1 0 624 0 1 18960
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_49
timestamp 1723858470
transform -1 0 624 0 -1 18960
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_50
timestamp 1723858470
transform -1 0 624 0 1 18170
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_51
timestamp 1723858470
transform -1 0 624 0 -1 18170
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_52
timestamp 1723858470
transform -1 0 624 0 1 17380
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_53
timestamp 1723858470
transform -1 0 624 0 -1 17380
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_54
timestamp 1723858470
transform -1 0 624 0 1 16590
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_55
timestamp 1723858470
transform -1 0 624 0 -1 16590
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_56
timestamp 1723858470
transform -1 0 624 0 1 15800
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_57
timestamp 1723858470
transform -1 0 624 0 -1 15800
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_58
timestamp 1723858470
transform -1 0 624 0 1 15010
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_59
timestamp 1723858470
transform -1 0 624 0 -1 15010
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_60
timestamp 1723858470
transform -1 0 624 0 1 14220
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_61
timestamp 1723858470
transform -1 0 624 0 -1 14220
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_62
timestamp 1723858470
transform -1 0 624 0 1 13430
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_63
timestamp 1723858470
transform -1 0 624 0 -1 13430
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_64
timestamp 1723858470
transform -1 0 624 0 1 26860
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_65
timestamp 1723858470
transform -1 0 624 0 -1 26860
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_66
timestamp 1723858470
transform -1 0 624 0 1 28440
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_67
timestamp 1723858470
transform -1 0 624 0 -1 28440
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_68
timestamp 1723858470
transform -1 0 624 0 1 27650
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_69
timestamp 1723858470
transform -1 0 624 0 -1 27650
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_70
timestamp 1723858470
transform -1 0 624 0 -1 38710
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_71
timestamp 1723858470
transform -1 0 624 0 1 37920
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_72
timestamp 1723858470
transform -1 0 624 0 -1 37920
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_73
timestamp 1723858470
transform -1 0 624 0 1 37130
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_74
timestamp 1723858470
transform -1 0 624 0 -1 37130
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_75
timestamp 1723858470
transform -1 0 624 0 1 36340
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_76
timestamp 1723858470
transform -1 0 624 0 -1 36340
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_77
timestamp 1723858470
transform -1 0 624 0 1 35550
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_78
timestamp 1723858470
transform -1 0 624 0 -1 35550
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_79
timestamp 1723858470
transform -1 0 624 0 1 34760
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_80
timestamp 1723858470
transform -1 0 624 0 -1 34760
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_81
timestamp 1723858470
transform -1 0 624 0 1 33970
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_82
timestamp 1723858470
transform -1 0 624 0 -1 33970
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_83
timestamp 1723858470
transform -1 0 624 0 1 33180
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_84
timestamp 1723858470
transform -1 0 624 0 -1 33180
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_85
timestamp 1723858470
transform -1 0 624 0 1 32390
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_86
timestamp 1723858470
transform -1 0 624 0 -1 32390
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_87
timestamp 1723858470
transform -1 0 624 0 1 31600
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_88
timestamp 1723858470
transform -1 0 624 0 -1 31600
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_89
timestamp 1723858470
transform -1 0 624 0 1 30810
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_90
timestamp 1723858470
transform -1 0 624 0 -1 30810
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_91
timestamp 1723858470
transform -1 0 624 0 1 30020
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_92
timestamp 1723858470
transform -1 0 624 0 -1 30020
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_93
timestamp 1723858470
transform -1 0 624 0 1 29230
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_94
timestamp 1723858470
transform -1 0 624 0 -1 29230
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_95
timestamp 1723858470
transform -1 0 624 0 -1 39500
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_96
timestamp 1723858470
transform -1 0 624 0 1 51350
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_97
timestamp 1723858470
transform -1 0 624 0 -1 51350
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_98
timestamp 1723858470
transform -1 0 624 0 1 50560
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_99
timestamp 1723858470
transform -1 0 624 0 -1 50560
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_100
timestamp 1723858470
transform -1 0 624 0 1 49770
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_101
timestamp 1723858470
transform -1 0 624 0 -1 49770
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_102
timestamp 1723858470
transform -1 0 624 0 1 48980
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_103
timestamp 1723858470
transform -1 0 624 0 -1 48980
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_104
timestamp 1723858470
transform -1 0 624 0 1 48190
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_105
timestamp 1723858470
transform -1 0 624 0 -1 48190
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_106
timestamp 1723858470
transform -1 0 624 0 1 47400
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_107
timestamp 1723858470
transform -1 0 624 0 -1 47400
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_108
timestamp 1723858470
transform -1 0 624 0 1 46610
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_109
timestamp 1723858470
transform -1 0 624 0 -1 46610
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_110
timestamp 1723858470
transform -1 0 624 0 1 45820
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_111
timestamp 1723858470
transform -1 0 624 0 -1 45820
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_112
timestamp 1723858470
transform -1 0 624 0 1 45030
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_113
timestamp 1723858470
transform -1 0 624 0 -1 45030
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_114
timestamp 1723858470
transform -1 0 624 0 1 44240
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_115
timestamp 1723858470
transform -1 0 624 0 -1 44240
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_116
timestamp 1723858470
transform -1 0 624 0 1 43450
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_117
timestamp 1723858470
transform -1 0 624 0 -1 43450
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_118
timestamp 1723858470
transform -1 0 624 0 1 42660
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_119
timestamp 1723858470
transform -1 0 624 0 -1 42660
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_120
timestamp 1723858470
transform -1 0 624 0 1 41870
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_121
timestamp 1723858470
transform -1 0 624 0 -1 41870
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_122
timestamp 1723858470
transform -1 0 624 0 1 41080
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_123
timestamp 1723858470
transform -1 0 624 0 -1 41080
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_124
timestamp 1723858470
transform -1 0 624 0 1 40290
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_125
timestamp 1723858470
transform -1 0 624 0 -1 40290
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_126
timestamp 1723858470
transform -1 0 624 0 1 39500
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_127
timestamp 1723858470
transform -1 0 624 0 1 38710
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_128
timestamp 1723858470
transform -1 0 624 0 1 26070
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_1  sky130_fd_bd_sram__openram_dp_cell_cap_row_129
timestamp 1723858470
transform -1 0 624 0 -1 26070
box -42 -55 624 371
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_0
timestamp 1723858470
transform 1 0 351 0 1 12840
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_1
timestamp 1723858470
transform 1 0 351 0 1 12603
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_2
timestamp 1723858470
transform 1 0 351 0 1 12366
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_3
timestamp 1723858470
transform 1 0 351 0 1 12050
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_4
timestamp 1723858470
transform 1 0 351 0 1 11813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_5
timestamp 1723858470
transform 1 0 351 0 1 11576
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_6
timestamp 1723858470
transform 1 0 351 0 1 11260
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_7
timestamp 1723858470
transform 1 0 351 0 1 11023
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_8
timestamp 1723858470
transform 1 0 351 0 1 10786
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_9
timestamp 1723858470
transform 1 0 351 0 1 10470
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_10
timestamp 1723858470
transform 1 0 351 0 1 10233
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_11
timestamp 1723858470
transform 1 0 351 0 1 9996
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_12
timestamp 1723858470
transform 1 0 351 0 1 9680
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_13
timestamp 1723858470
transform 1 0 351 0 1 9443
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_14
timestamp 1723858470
transform 1 0 351 0 1 9206
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_15
timestamp 1723858470
transform 1 0 351 0 1 8890
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_16
timestamp 1723858470
transform 1 0 351 0 1 8653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_17
timestamp 1723858470
transform 1 0 351 0 1 8416
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_18
timestamp 1723858470
transform 1 0 351 0 1 8100
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_19
timestamp 1723858470
transform 1 0 351 0 1 7863
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_20
timestamp 1723858470
transform 1 0 351 0 1 7626
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_21
timestamp 1723858470
transform 1 0 351 0 1 7310
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_22
timestamp 1723858470
transform 1 0 351 0 1 7073
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_23
timestamp 1723858470
transform 1 0 351 0 1 6836
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_24
timestamp 1723858470
transform 1 0 351 0 1 6520
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_25
timestamp 1723858470
transform 1 0 351 0 1 6283
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_26
timestamp 1723858470
transform 1 0 351 0 1 6046
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_27
timestamp 1723858470
transform 1 0 351 0 1 5730
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_28
timestamp 1723858470
transform 1 0 351 0 1 5493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_29
timestamp 1723858470
transform 1 0 351 0 1 5256
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_30
timestamp 1723858470
transform 1 0 351 0 1 4940
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_31
timestamp 1723858470
transform 1 0 351 0 1 4703
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_32
timestamp 1723858470
transform 1 0 351 0 1 4466
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_33
timestamp 1723858470
transform 1 0 351 0 1 4150
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_34
timestamp 1723858470
transform 1 0 351 0 1 3913
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_35
timestamp 1723858470
transform 1 0 351 0 1 3676
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_36
timestamp 1723858470
transform 1 0 351 0 1 3360
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_37
timestamp 1723858470
transform 1 0 351 0 1 3123
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_38
timestamp 1723858470
transform 1 0 351 0 1 2886
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_39
timestamp 1723858470
transform 1 0 351 0 1 2570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_40
timestamp 1723858470
transform 1 0 351 0 1 2333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_41
timestamp 1723858470
transform 1 0 351 0 1 2096
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_42
timestamp 1723858470
transform 1 0 351 0 1 1780
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_43
timestamp 1723858470
transform 1 0 351 0 1 1543
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_44
timestamp 1723858470
transform 1 0 351 0 1 1306
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_45
timestamp 1723858470
transform 1 0 351 0 1 753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_46
timestamp 1723858470
transform 1 0 351 0 1 990
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_47
timestamp 1723858470
transform 1 0 351 0 1 13630
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_48
timestamp 1723858470
transform 1 0 351 0 1 13946
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_49
timestamp 1723858470
transform 1 0 351 0 1 13393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_50
timestamp 1723858470
transform 1 0 351 0 1 25796
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_51
timestamp 1723858470
transform 1 0 351 0 1 25480
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_52
timestamp 1723858470
transform 1 0 351 0 1 25243
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_53
timestamp 1723858470
transform 1 0 351 0 1 25006
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_54
timestamp 1723858470
transform 1 0 351 0 1 24690
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_55
timestamp 1723858470
transform 1 0 351 0 1 24453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_56
timestamp 1723858470
transform 1 0 351 0 1 24216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_57
timestamp 1723858470
transform 1 0 351 0 1 23900
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_58
timestamp 1723858470
transform 1 0 351 0 1 23663
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_59
timestamp 1723858470
transform 1 0 351 0 1 23426
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_60
timestamp 1723858470
transform 1 0 351 0 1 23110
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_61
timestamp 1723858470
transform 1 0 351 0 1 22873
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_62
timestamp 1723858470
transform 1 0 351 0 1 22636
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_63
timestamp 1723858470
transform 1 0 351 0 1 22320
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_64
timestamp 1723858470
transform 1 0 351 0 1 22083
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_65
timestamp 1723858470
transform 1 0 351 0 1 21846
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_66
timestamp 1723858470
transform 1 0 351 0 1 21530
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_67
timestamp 1723858470
transform 1 0 351 0 1 21293
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_68
timestamp 1723858470
transform 1 0 351 0 1 21056
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_69
timestamp 1723858470
transform 1 0 351 0 1 20740
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_70
timestamp 1723858470
transform 1 0 351 0 1 20503
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_71
timestamp 1723858470
transform 1 0 351 0 1 20266
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_72
timestamp 1723858470
transform 1 0 351 0 1 19950
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_73
timestamp 1723858470
transform 1 0 351 0 1 19713
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_74
timestamp 1723858470
transform 1 0 351 0 1 19476
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_75
timestamp 1723858470
transform 1 0 351 0 1 19160
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_76
timestamp 1723858470
transform 1 0 351 0 1 18923
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_77
timestamp 1723858470
transform 1 0 351 0 1 18686
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_78
timestamp 1723858470
transform 1 0 351 0 1 18370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_79
timestamp 1723858470
transform 1 0 351 0 1 18133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_80
timestamp 1723858470
transform 1 0 351 0 1 17896
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_81
timestamp 1723858470
transform 1 0 351 0 1 17580
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_82
timestamp 1723858470
transform 1 0 351 0 1 17343
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_83
timestamp 1723858470
transform 1 0 351 0 1 17106
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_84
timestamp 1723858470
transform 1 0 351 0 1 16790
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_85
timestamp 1723858470
transform 1 0 351 0 1 16553
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_86
timestamp 1723858470
transform 1 0 351 0 1 16316
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_87
timestamp 1723858470
transform 1 0 351 0 1 16000
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_88
timestamp 1723858470
transform 1 0 351 0 1 15763
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_89
timestamp 1723858470
transform 1 0 351 0 1 15526
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_90
timestamp 1723858470
transform 1 0 351 0 1 15210
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_91
timestamp 1723858470
transform 1 0 351 0 1 14973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_92
timestamp 1723858470
transform 1 0 351 0 1 14736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_93
timestamp 1723858470
transform 1 0 351 0 1 14420
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_94
timestamp 1723858470
transform 1 0 351 0 1 14183
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_95
timestamp 1723858470
transform 1 0 351 0 1 13156
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_96
timestamp 1723858470
transform 1 0 351 0 1 32590
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_97
timestamp 1723858470
transform 1 0 351 0 1 32116
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_98
timestamp 1723858470
transform 1 0 351 0 1 31800
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_99
timestamp 1723858470
transform 1 0 351 0 1 31563
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_100
timestamp 1723858470
transform 1 0 351 0 1 31326
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_101
timestamp 1723858470
transform 1 0 351 0 1 31010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_102
timestamp 1723858470
transform 1 0 351 0 1 30773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_103
timestamp 1723858470
transform 1 0 351 0 1 30536
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_104
timestamp 1723858470
transform 1 0 351 0 1 30220
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_105
timestamp 1723858470
transform 1 0 351 0 1 29983
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_106
timestamp 1723858470
transform 1 0 351 0 1 29746
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_107
timestamp 1723858470
transform 1 0 351 0 1 29430
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_108
timestamp 1723858470
transform 1 0 351 0 1 29193
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_109
timestamp 1723858470
transform 1 0 351 0 1 28956
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_110
timestamp 1723858470
transform 1 0 351 0 1 28640
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_111
timestamp 1723858470
transform 1 0 351 0 1 28403
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_112
timestamp 1723858470
transform 1 0 351 0 1 28166
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_113
timestamp 1723858470
transform 1 0 351 0 1 27850
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_114
timestamp 1723858470
transform 1 0 351 0 1 27613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_115
timestamp 1723858470
transform 1 0 351 0 1 27376
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_116
timestamp 1723858470
transform 1 0 351 0 1 27060
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_117
timestamp 1723858470
transform 1 0 351 0 1 26823
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_118
timestamp 1723858470
transform 1 0 351 0 1 26586
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_119
timestamp 1723858470
transform 1 0 351 0 1 26270
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_120
timestamp 1723858470
transform 1 0 351 0 1 38673
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_121
timestamp 1723858470
transform 1 0 351 0 1 38436
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_122
timestamp 1723858470
transform 1 0 351 0 1 38120
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_123
timestamp 1723858470
transform 1 0 351 0 1 37883
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_124
timestamp 1723858470
transform 1 0 351 0 1 37646
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_125
timestamp 1723858470
transform 1 0 351 0 1 37330
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_126
timestamp 1723858470
transform 1 0 351 0 1 37093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_127
timestamp 1723858470
transform 1 0 351 0 1 36856
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_128
timestamp 1723858470
transform 1 0 351 0 1 36540
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_129
timestamp 1723858470
transform 1 0 351 0 1 36303
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_130
timestamp 1723858470
transform 1 0 351 0 1 36066
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_131
timestamp 1723858470
transform 1 0 351 0 1 35750
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_132
timestamp 1723858470
transform 1 0 351 0 1 35513
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_133
timestamp 1723858470
transform 1 0 351 0 1 35276
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_134
timestamp 1723858470
transform 1 0 351 0 1 34960
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_135
timestamp 1723858470
transform 1 0 351 0 1 34723
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_136
timestamp 1723858470
transform 1 0 351 0 1 34486
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_137
timestamp 1723858470
transform 1 0 351 0 1 34170
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_138
timestamp 1723858470
transform 1 0 351 0 1 33933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_139
timestamp 1723858470
transform 1 0 351 0 1 33696
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_140
timestamp 1723858470
transform 1 0 351 0 1 33380
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_141
timestamp 1723858470
transform 1 0 351 0 1 33143
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_142
timestamp 1723858470
transform 1 0 351 0 1 32906
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_143
timestamp 1723858470
transform 1 0 351 0 1 32353
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_144
timestamp 1723858470
transform 1 0 351 0 1 51313
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_145
timestamp 1723858470
transform 1 0 351 0 1 51076
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_146
timestamp 1723858470
transform 1 0 351 0 1 50760
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_147
timestamp 1723858470
transform 1 0 351 0 1 50523
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_148
timestamp 1723858470
transform 1 0 351 0 1 50286
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_149
timestamp 1723858470
transform 1 0 351 0 1 49970
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_150
timestamp 1723858470
transform 1 0 351 0 1 49733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_151
timestamp 1723858470
transform 1 0 351 0 1 49496
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_152
timestamp 1723858470
transform 1 0 351 0 1 49180
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_153
timestamp 1723858470
transform 1 0 351 0 1 48943
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_154
timestamp 1723858470
transform 1 0 351 0 1 48706
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_155
timestamp 1723858470
transform 1 0 351 0 1 48390
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_156
timestamp 1723858470
transform 1 0 351 0 1 48153
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_157
timestamp 1723858470
transform 1 0 351 0 1 47916
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_158
timestamp 1723858470
transform 1 0 351 0 1 47600
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_159
timestamp 1723858470
transform 1 0 351 0 1 47363
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_160
timestamp 1723858470
transform 1 0 351 0 1 47126
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_161
timestamp 1723858470
transform 1 0 351 0 1 46810
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_162
timestamp 1723858470
transform 1 0 351 0 1 46573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_163
timestamp 1723858470
transform 1 0 351 0 1 46336
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_164
timestamp 1723858470
transform 1 0 351 0 1 46020
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_165
timestamp 1723858470
transform 1 0 351 0 1 45783
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_166
timestamp 1723858470
transform 1 0 351 0 1 45546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_167
timestamp 1723858470
transform 1 0 351 0 1 45230
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_168
timestamp 1723858470
transform 1 0 351 0 1 44993
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_169
timestamp 1723858470
transform 1 0 351 0 1 44756
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_170
timestamp 1723858470
transform 1 0 351 0 1 44440
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_171
timestamp 1723858470
transform 1 0 351 0 1 44203
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_172
timestamp 1723858470
transform 1 0 351 0 1 43966
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_173
timestamp 1723858470
transform 1 0 351 0 1 43650
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_174
timestamp 1723858470
transform 1 0 351 0 1 43413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_175
timestamp 1723858470
transform 1 0 351 0 1 43176
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_176
timestamp 1723858470
transform 1 0 351 0 1 42860
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_177
timestamp 1723858470
transform 1 0 351 0 1 42623
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_178
timestamp 1723858470
transform 1 0 351 0 1 42386
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_179
timestamp 1723858470
transform 1 0 351 0 1 42070
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_180
timestamp 1723858470
transform 1 0 351 0 1 41833
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_181
timestamp 1723858470
transform 1 0 351 0 1 41596
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_182
timestamp 1723858470
transform 1 0 351 0 1 41280
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_183
timestamp 1723858470
transform 1 0 351 0 1 41043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_184
timestamp 1723858470
transform 1 0 351 0 1 40806
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_185
timestamp 1723858470
transform 1 0 351 0 1 40490
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_186
timestamp 1723858470
transform 1 0 351 0 1 40253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_187
timestamp 1723858470
transform 1 0 351 0 1 40016
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_188
timestamp 1723858470
transform 1 0 351 0 1 39700
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_189
timestamp 1723858470
transform 1 0 351 0 1 39463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_190
timestamp 1723858470
transform 1 0 351 0 1 39226
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_191
timestamp 1723858470
transform 1 0 351 0 1 38910
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_192
timestamp 1723858470
transform 1 0 351 0 1 26033
box 0 0 1 1
<< labels >>
rlabel metal3 s 335 29418 433 29516 4 gnd
port 1 nsew
rlabel metal3 s 335 47351 433 47449 4 gnd
port 1 nsew
rlabel metal3 s 335 35738 433 35836 4 gnd
port 1 nsew
rlabel metal3 s 335 44744 433 44842 4 gnd
port 1 nsew
rlabel metal3 s 335 39451 433 39549 4 gnd
port 1 nsew
rlabel metal3 s 335 28628 433 28726 4 gnd
port 1 nsew
rlabel metal3 s 335 48141 433 48239 4 gnd
port 1 nsew
rlabel metal3 s 335 34711 433 34809 4 gnd
port 1 nsew
rlabel metal3 s 335 35501 433 35599 4 gnd
port 1 nsew
rlabel metal3 s 335 34948 433 35046 4 gnd
port 1 nsew
rlabel metal3 s 335 45771 433 45869 4 gnd
port 1 nsew
rlabel metal3 s 335 40794 433 40892 4 gnd
port 1 nsew
rlabel metal3 s 335 47904 433 48002 4 gnd
port 1 nsew
rlabel metal3 s 335 38661 433 38759 4 gnd
port 1 nsew
rlabel metal3 s 335 44981 433 45079 4 gnd
port 1 nsew
rlabel metal3 s 335 26811 433 26909 4 gnd
port 1 nsew
rlabel metal3 s 335 26258 433 26356 4 gnd
port 1 nsew
rlabel metal3 s 335 36528 433 36626 4 gnd
port 1 nsew
rlabel metal3 s 335 49484 433 49582 4 gnd
port 1 nsew
rlabel metal3 s 335 27601 433 27699 4 gnd
port 1 nsew
rlabel metal3 s 335 39688 433 39786 4 gnd
port 1 nsew
rlabel metal3 s 335 32894 433 32992 4 gnd
port 1 nsew
rlabel metal3 s 335 27364 433 27462 4 gnd
port 1 nsew
rlabel metal3 s 335 31788 433 31886 4 gnd
port 1 nsew
rlabel metal3 s 335 50274 433 50372 4 gnd
port 1 nsew
rlabel metal3 s 335 44428 433 44526 4 gnd
port 1 nsew
rlabel metal3 s 335 33131 433 33229 4 gnd
port 1 nsew
rlabel metal3 s 335 43401 433 43499 4 gnd
port 1 nsew
rlabel metal3 s 335 41268 433 41366 4 gnd
port 1 nsew
rlabel metal3 s 335 40478 433 40576 4 gnd
port 1 nsew
rlabel metal3 s 335 33684 433 33782 4 gnd
port 1 nsew
rlabel metal3 s 335 37871 433 37969 4 gnd
port 1 nsew
rlabel metal3 s 335 43164 433 43262 4 gnd
port 1 nsew
rlabel metal3 s 335 28154 433 28252 4 gnd
port 1 nsew
rlabel metal3 s 335 30761 433 30859 4 gnd
port 1 nsew
rlabel metal3 s 335 50748 433 50846 4 gnd
port 1 nsew
rlabel metal3 s 335 33368 433 33466 4 gnd
port 1 nsew
rlabel metal3 s 335 36291 433 36389 4 gnd
port 1 nsew
rlabel metal3 s 335 46561 433 46659 4 gnd
port 1 nsew
rlabel metal3 s 335 42374 433 42472 4 gnd
port 1 nsew
rlabel metal3 s 335 29971 433 30069 4 gnd
port 1 nsew
rlabel metal3 s 335 46324 433 46422 4 gnd
port 1 nsew
rlabel metal3 s 335 42058 433 42156 4 gnd
port 1 nsew
rlabel metal3 s 335 37081 433 37179 4 gnd
port 1 nsew
rlabel metal3 s 335 51064 433 51162 4 gnd
port 1 nsew
rlabel metal3 s 335 34474 433 34572 4 gnd
port 1 nsew
rlabel metal3 s 335 31314 433 31412 4 gnd
port 1 nsew
rlabel metal3 s 335 28391 433 28489 4 gnd
port 1 nsew
rlabel metal3 s 335 39214 433 39312 4 gnd
port 1 nsew
rlabel metal3 s 335 44191 433 44289 4 gnd
port 1 nsew
rlabel metal3 s 335 49958 433 50056 4 gnd
port 1 nsew
rlabel metal3 s 335 30524 433 30622 4 gnd
port 1 nsew
rlabel metal3 s 335 48378 433 48476 4 gnd
port 1 nsew
rlabel metal3 s 335 30208 433 30306 4 gnd
port 1 nsew
rlabel metal3 s 335 48694 433 48792 4 gnd
port 1 nsew
rlabel metal3 s 335 33921 433 34019 4 gnd
port 1 nsew
rlabel metal3 s 335 41584 433 41682 4 gnd
port 1 nsew
rlabel metal3 s 335 46008 433 46106 4 gnd
port 1 nsew
rlabel metal3 s 335 48931 433 49029 4 gnd
port 1 nsew
rlabel metal3 s 335 51301 433 51399 4 gnd
port 1 nsew
rlabel metal3 s 335 38898 433 38996 4 gnd
port 1 nsew
rlabel metal3 s 335 31551 433 31649 4 gnd
port 1 nsew
rlabel metal3 s 335 26574 433 26672 4 gnd
port 1 nsew
rlabel metal3 s 335 30998 433 31096 4 gnd
port 1 nsew
rlabel metal3 s 335 37318 433 37416 4 gnd
port 1 nsew
rlabel metal3 s 335 27048 433 27146 4 gnd
port 1 nsew
rlabel metal3 s 335 40241 433 40339 4 gnd
port 1 nsew
rlabel metal3 s 335 32104 433 32202 4 gnd
port 1 nsew
rlabel metal3 s 335 40004 433 40102 4 gnd
port 1 nsew
rlabel metal3 s 335 46798 433 46896 4 gnd
port 1 nsew
rlabel metal3 s 335 41821 433 41919 4 gnd
port 1 nsew
rlabel metal3 s 335 49721 433 49819 4 gnd
port 1 nsew
rlabel metal3 s 335 36054 433 36152 4 gnd
port 1 nsew
rlabel metal3 s 335 49168 433 49266 4 gnd
port 1 nsew
rlabel metal3 s 335 32341 433 32439 4 gnd
port 1 nsew
rlabel metal3 s 335 38108 433 38206 4 gnd
port 1 nsew
rlabel metal3 s 335 43954 433 44052 4 gnd
port 1 nsew
rlabel metal3 s 335 28944 433 29042 4 gnd
port 1 nsew
rlabel metal3 s 335 43638 433 43736 4 gnd
port 1 nsew
rlabel metal3 s 335 36844 433 36942 4 gnd
port 1 nsew
rlabel metal3 s 335 50511 433 50609 4 gnd
port 1 nsew
rlabel metal3 s 335 32578 433 32676 4 gnd
port 1 nsew
rlabel metal3 s 335 27838 433 27936 4 gnd
port 1 nsew
rlabel metal3 s 335 45218 433 45316 4 gnd
port 1 nsew
rlabel metal3 s 335 35264 433 35362 4 gnd
port 1 nsew
rlabel metal3 s 335 47588 433 47686 4 gnd
port 1 nsew
rlabel metal3 s 335 47114 433 47212 4 gnd
port 1 nsew
rlabel metal3 s 335 34158 433 34256 4 gnd
port 1 nsew
rlabel metal3 s 335 41031 433 41129 4 gnd
port 1 nsew
rlabel metal3 s 335 42848 433 42946 4 gnd
port 1 nsew
rlabel metal3 s 335 37634 433 37732 4 gnd
port 1 nsew
rlabel metal3 s 335 29181 433 29279 4 gnd
port 1 nsew
rlabel metal3 s 335 38424 433 38522 4 gnd
port 1 nsew
rlabel metal3 s 335 45534 433 45632 4 gnd
port 1 nsew
rlabel metal3 s 335 42611 433 42709 4 gnd
port 1 nsew
rlabel metal3 s 335 29734 433 29832 4 gnd
port 1 nsew
rlabel metal3 s 335 19701 433 19799 4 gnd
port 1 nsew
rlabel metal3 s 335 1531 433 1629 4 gnd
port 1 nsew
rlabel metal3 s 335 21518 433 21616 4 gnd
port 1 nsew
rlabel metal3 s 335 24994 433 25092 4 gnd
port 1 nsew
rlabel metal3 s 335 10221 433 10319 4 gnd
port 1 nsew
rlabel metal3 s 335 18911 433 19009 4 gnd
port 1 nsew
rlabel metal3 s 335 16778 433 16876 4 gnd
port 1 nsew
rlabel metal3 s 335 15751 433 15849 4 gnd
port 1 nsew
rlabel metal3 s 335 4928 433 5026 4 gnd
port 1 nsew
rlabel metal3 s 335 16304 433 16402 4 gnd
port 1 nsew
rlabel metal3 s 335 19464 433 19562 4 gnd
port 1 nsew
rlabel metal3 s 335 22071 433 22169 4 gnd
port 1 nsew
rlabel metal3 s 335 12828 433 12926 4 gnd
port 1 nsew
rlabel metal3 s 335 14961 433 15059 4 gnd
port 1 nsew
rlabel metal3 s 335 12591 433 12689 4 gnd
port 1 nsew
rlabel metal3 s 335 4691 433 4789 4 gnd
port 1 nsew
rlabel metal3 s 335 2874 433 2972 4 gnd
port 1 nsew
rlabel metal3 s 335 18674 433 18772 4 gnd
port 1 nsew
rlabel metal3 s 335 25784 433 25882 4 gnd
port 1 nsew
rlabel metal3 s 335 741 433 839 4 gnd
port 1 nsew
rlabel metal3 s 335 7298 433 7396 4 gnd
port 1 nsew
rlabel metal3 s 335 4454 433 4552 4 gnd
port 1 nsew
rlabel metal3 s 335 9668 433 9766 4 gnd
port 1 nsew
rlabel metal3 s 335 11011 433 11109 4 gnd
port 1 nsew
rlabel metal3 s 335 5481 433 5579 4 gnd
port 1 nsew
rlabel metal3 s 335 13381 433 13479 4 gnd
port 1 nsew
rlabel metal3 s 335 23414 433 23512 4 gnd
port 1 nsew
rlabel metal3 s 335 17094 433 17192 4 gnd
port 1 nsew
rlabel metal3 s 335 2084 433 2182 4 gnd
port 1 nsew
rlabel metal3 s 335 24441 433 24539 4 gnd
port 1 nsew
rlabel metal3 s 335 14408 433 14506 4 gnd
port 1 nsew
rlabel metal3 s 335 19938 433 20036 4 gnd
port 1 nsew
rlabel metal3 s 335 16541 433 16639 4 gnd
port 1 nsew
rlabel metal3 s 335 14171 433 14269 4 gnd
port 1 nsew
rlabel metal3 s 335 20254 433 20352 4 gnd
port 1 nsew
rlabel metal3 s 335 7061 433 7159 4 gnd
port 1 nsew
rlabel metal3 s 335 2321 433 2419 4 gnd
port 1 nsew
rlabel metal3 s 335 18121 433 18219 4 gnd
port 1 nsew
rlabel metal3 s 335 22624 433 22722 4 gnd
port 1 nsew
rlabel metal3 s 335 11801 433 11899 4 gnd
port 1 nsew
rlabel metal3 s 335 17331 433 17429 4 gnd
port 1 nsew
rlabel metal3 s 335 3664 433 3762 4 gnd
port 1 nsew
rlabel metal3 s 335 10458 433 10556 4 gnd
port 1 nsew
rlabel metal3 s 335 23651 433 23749 4 gnd
port 1 nsew
rlabel metal3 s 335 10774 433 10872 4 gnd
port 1 nsew
rlabel metal3 s 335 9194 433 9292 4 gnd
port 1 nsew
rlabel metal3 s 335 9984 433 10082 4 gnd
port 1 nsew
rlabel metal3 s 335 3111 433 3209 4 gnd
port 1 nsew
rlabel metal3 s 335 6271 433 6369 4 gnd
port 1 nsew
rlabel metal3 s 335 5718 433 5816 4 gnd
port 1 nsew
rlabel metal3 s 335 22861 433 22959 4 gnd
port 1 nsew
rlabel metal3 s 335 15514 433 15612 4 gnd
port 1 nsew
rlabel metal3 s 335 6034 433 6132 4 gnd
port 1 nsew
rlabel metal3 s 335 22308 433 22406 4 gnd
port 1 nsew
rlabel metal3 s 335 2558 433 2656 4 gnd
port 1 nsew
rlabel metal3 s 335 12354 433 12452 4 gnd
port 1 nsew
rlabel metal3 s 335 20728 433 20826 4 gnd
port 1 nsew
rlabel metal3 s 335 13618 433 13716 4 gnd
port 1 nsew
rlabel metal3 s 335 23098 433 23196 4 gnd
port 1 nsew
rlabel metal3 s 335 8878 433 8976 4 gnd
port 1 nsew
rlabel metal3 s 335 1768 433 1866 4 gnd
port 1 nsew
rlabel metal3 s 335 8641 433 8739 4 gnd
port 1 nsew
rlabel metal3 s 335 17884 433 17982 4 gnd
port 1 nsew
rlabel metal3 s 335 21044 433 21142 4 gnd
port 1 nsew
rlabel metal3 s 335 23888 433 23986 4 gnd
port 1 nsew
rlabel metal3 s 335 1294 433 1392 4 gnd
port 1 nsew
rlabel metal3 s 335 13934 433 14032 4 gnd
port 1 nsew
rlabel metal3 s 335 21834 433 21932 4 gnd
port 1 nsew
rlabel metal3 s 335 13144 433 13242 4 gnd
port 1 nsew
rlabel metal3 s 335 9431 433 9529 4 gnd
port 1 nsew
rlabel metal3 s 335 15988 433 16086 4 gnd
port 1 nsew
rlabel metal3 s 335 26021 433 26119 4 gnd
port 1 nsew
rlabel metal3 s 335 18358 433 18456 4 gnd
port 1 nsew
rlabel metal3 s 335 6824 433 6922 4 gnd
port 1 nsew
rlabel metal3 s 335 14724 433 14822 4 gnd
port 1 nsew
rlabel metal3 s 335 25468 433 25566 4 gnd
port 1 nsew
rlabel metal3 s 335 7614 433 7712 4 gnd
port 1 nsew
rlabel metal3 s 335 8404 433 8502 4 gnd
port 1 nsew
rlabel metal3 s 335 25231 433 25329 4 gnd
port 1 nsew
rlabel metal3 s 335 3901 433 3999 4 gnd
port 1 nsew
rlabel metal3 s 335 17568 433 17666 4 gnd
port 1 nsew
rlabel metal3 s 335 978 433 1076 4 gnd
port 1 nsew
rlabel metal3 s 335 19148 433 19246 4 gnd
port 1 nsew
rlabel metal3 s 335 11248 433 11346 4 gnd
port 1 nsew
rlabel metal3 s 335 11564 433 11662 4 gnd
port 1 nsew
rlabel metal3 s 335 24678 433 24776 4 gnd
port 1 nsew
rlabel metal3 s 335 24204 433 24302 4 gnd
port 1 nsew
rlabel metal3 s 335 5244 433 5342 4 gnd
port 1 nsew
rlabel metal3 s 335 12038 433 12136 4 gnd
port 1 nsew
rlabel metal3 s 335 20491 433 20589 4 gnd
port 1 nsew
rlabel metal3 s 335 7851 433 7949 4 gnd
port 1 nsew
rlabel metal3 s 335 15198 433 15296 4 gnd
port 1 nsew
rlabel metal3 s 335 6508 433 6606 4 gnd
port 1 nsew
rlabel metal3 s 335 21281 433 21379 4 gnd
port 1 nsew
rlabel metal3 s 335 3348 433 3446 4 gnd
port 1 nsew
rlabel metal3 s 335 4138 433 4236 4 gnd
port 1 nsew
rlabel metal3 s 335 8088 433 8186 4 gnd
port 1 nsew
rlabel metal2 s 0 39033 28 39081 4 wl0_97
port 2 nsew
rlabel metal2 s 0 38813 28 38861 4 wl1_97
port 3 nsew
rlabel metal2 s 0 39129 28 39177 4 wl0_98
port 4 nsew
rlabel metal2 s 0 39349 28 39397 4 wl1_98
port 5 nsew
rlabel metal2 s 0 39823 28 39871 4 wl0_99
port 6 nsew
rlabel metal2 s 0 39603 28 39651 4 wl1_99
port 7 nsew
rlabel metal2 s 0 39919 28 39967 4 wl0_100
port 8 nsew
rlabel metal2 s 0 40139 28 40187 4 wl1_100
port 9 nsew
rlabel metal2 s 0 40613 28 40661 4 wl0_101
port 10 nsew
rlabel metal2 s 0 40393 28 40441 4 wl1_101
port 11 nsew
rlabel metal2 s 0 40709 28 40757 4 wl0_102
port 12 nsew
rlabel metal2 s 0 40929 28 40977 4 wl1_102
port 13 nsew
rlabel metal2 s 0 41403 28 41451 4 wl0_103
port 14 nsew
rlabel metal2 s 0 41183 28 41231 4 wl1_103
port 15 nsew
rlabel metal2 s 0 41499 28 41547 4 wl0_104
port 16 nsew
rlabel metal2 s 0 41719 28 41767 4 wl1_104
port 17 nsew
rlabel metal2 s 0 42193 28 42241 4 wl0_105
port 18 nsew
rlabel metal2 s 0 41973 28 42021 4 wl1_105
port 19 nsew
rlabel metal2 s 0 42289 28 42337 4 wl0_106
port 20 nsew
rlabel metal2 s 0 42509 28 42557 4 wl1_106
port 21 nsew
rlabel metal2 s 0 42983 28 43031 4 wl0_107
port 22 nsew
rlabel metal2 s 0 42763 28 42811 4 wl1_107
port 23 nsew
rlabel metal2 s 0 43079 28 43127 4 wl0_108
port 24 nsew
rlabel metal2 s 0 43299 28 43347 4 wl1_108
port 25 nsew
rlabel metal2 s 0 43773 28 43821 4 wl0_109
port 26 nsew
rlabel metal2 s 0 43553 28 43601 4 wl1_109
port 27 nsew
rlabel metal2 s 0 43869 28 43917 4 wl0_110
port 28 nsew
rlabel metal2 s 0 44089 28 44137 4 wl1_110
port 29 nsew
rlabel metal2 s 0 44563 28 44611 4 wl0_111
port 30 nsew
rlabel metal2 s 0 44343 28 44391 4 wl1_111
port 31 nsew
rlabel metal2 s 0 44659 28 44707 4 wl0_112
port 32 nsew
rlabel metal2 s 0 44879 28 44927 4 wl1_112
port 33 nsew
rlabel metal2 s 0 45353 28 45401 4 wl0_113
port 34 nsew
rlabel metal2 s 0 45133 28 45181 4 wl1_113
port 35 nsew
rlabel metal2 s 0 45449 28 45497 4 wl0_114
port 36 nsew
rlabel metal2 s 0 45669 28 45717 4 wl1_114
port 37 nsew
rlabel metal2 s 0 46143 28 46191 4 wl0_115
port 38 nsew
rlabel metal2 s 0 45923 28 45971 4 wl1_115
port 39 nsew
rlabel metal2 s 0 46239 28 46287 4 wl0_116
port 40 nsew
rlabel metal2 s 0 46459 28 46507 4 wl1_116
port 41 nsew
rlabel metal2 s 0 46933 28 46981 4 wl0_117
port 42 nsew
rlabel metal2 s 0 46713 28 46761 4 wl1_117
port 43 nsew
rlabel metal2 s 0 47029 28 47077 4 wl0_118
port 44 nsew
rlabel metal2 s 0 47249 28 47297 4 wl1_118
port 45 nsew
rlabel metal2 s 0 47723 28 47771 4 wl0_119
port 46 nsew
rlabel metal2 s 0 47503 28 47551 4 wl1_119
port 47 nsew
rlabel metal2 s 0 47819 28 47867 4 wl0_120
port 48 nsew
rlabel metal2 s 0 48039 28 48087 4 wl1_120
port 49 nsew
rlabel metal2 s 0 48513 28 48561 4 wl0_121
port 50 nsew
rlabel metal2 s 0 48293 28 48341 4 wl1_121
port 51 nsew
rlabel metal2 s 0 48609 28 48657 4 wl0_122
port 52 nsew
rlabel metal2 s 0 48829 28 48877 4 wl1_122
port 53 nsew
rlabel metal2 s 0 49303 28 49351 4 wl0_123
port 54 nsew
rlabel metal2 s 0 49083 28 49131 4 wl1_123
port 55 nsew
rlabel metal2 s 0 49399 28 49447 4 wl0_124
port 56 nsew
rlabel metal2 s 0 49619 28 49667 4 wl1_124
port 57 nsew
rlabel metal2 s 0 50093 28 50141 4 wl0_125
port 58 nsew
rlabel metal2 s 0 49873 28 49921 4 wl1_125
port 59 nsew
rlabel metal2 s 0 50189 28 50237 4 wl0_126
port 60 nsew
rlabel metal2 s 0 50409 28 50457 4 wl1_126
port 61 nsew
rlabel metal2 s 0 50883 28 50931 4 wl0_127
port 62 nsew
rlabel metal2 s 0 50663 28 50711 4 wl1_127
port 63 nsew
rlabel metal2 s 0 50979 28 51027 4 wl0_128
port 64 nsew
rlabel metal2 s 0 51199 28 51247 4 wl1_128
port 65 nsew
rlabel metal2 s 0 26393 28 26441 4 wl0_65
port 66 nsew
rlabel metal2 s 0 26173 28 26221 4 wl1_65
port 67 nsew
rlabel metal2 s 0 26489 28 26537 4 wl0_66
port 68 nsew
rlabel metal2 s 0 26709 28 26757 4 wl1_66
port 69 nsew
rlabel metal2 s 0 27183 28 27231 4 wl0_67
port 70 nsew
rlabel metal2 s 0 26963 28 27011 4 wl1_67
port 71 nsew
rlabel metal2 s 0 27279 28 27327 4 wl0_68
port 72 nsew
rlabel metal2 s 0 27499 28 27547 4 wl1_68
port 73 nsew
rlabel metal2 s 0 27973 28 28021 4 wl0_69
port 74 nsew
rlabel metal2 s 0 27753 28 27801 4 wl1_69
port 75 nsew
rlabel metal2 s 0 28069 28 28117 4 wl0_70
port 76 nsew
rlabel metal2 s 0 28289 28 28337 4 wl1_70
port 77 nsew
rlabel metal2 s 0 28763 28 28811 4 wl0_71
port 78 nsew
rlabel metal2 s 0 28543 28 28591 4 wl1_71
port 79 nsew
rlabel metal2 s 0 28859 28 28907 4 wl0_72
port 80 nsew
rlabel metal2 s 0 29079 28 29127 4 wl1_72
port 81 nsew
rlabel metal2 s 0 29553 28 29601 4 wl0_73
port 82 nsew
rlabel metal2 s 0 29333 28 29381 4 wl1_73
port 83 nsew
rlabel metal2 s 0 29649 28 29697 4 wl0_74
port 84 nsew
rlabel metal2 s 0 29869 28 29917 4 wl1_74
port 85 nsew
rlabel metal2 s 0 30343 28 30391 4 wl0_75
port 86 nsew
rlabel metal2 s 0 30123 28 30171 4 wl1_75
port 87 nsew
rlabel metal2 s 0 30439 28 30487 4 wl0_76
port 88 nsew
rlabel metal2 s 0 30659 28 30707 4 wl1_76
port 89 nsew
rlabel metal2 s 0 31133 28 31181 4 wl0_77
port 90 nsew
rlabel metal2 s 0 30913 28 30961 4 wl1_77
port 91 nsew
rlabel metal2 s 0 31229 28 31277 4 wl0_78
port 92 nsew
rlabel metal2 s 0 31449 28 31497 4 wl1_78
port 93 nsew
rlabel metal2 s 0 31923 28 31971 4 wl0_79
port 94 nsew
rlabel metal2 s 0 31703 28 31751 4 wl1_79
port 95 nsew
rlabel metal2 s 0 32019 28 32067 4 wl0_80
port 96 nsew
rlabel metal2 s 0 32239 28 32287 4 wl1_80
port 97 nsew
rlabel metal2 s 0 32713 28 32761 4 wl0_81
port 98 nsew
rlabel metal2 s 0 32493 28 32541 4 wl1_81
port 99 nsew
rlabel metal2 s 0 32809 28 32857 4 wl0_82
port 100 nsew
rlabel metal2 s 0 33029 28 33077 4 wl1_82
port 101 nsew
rlabel metal2 s 0 33503 28 33551 4 wl0_83
port 102 nsew
rlabel metal2 s 0 33283 28 33331 4 wl1_83
port 103 nsew
rlabel metal2 s 0 33599 28 33647 4 wl0_84
port 104 nsew
rlabel metal2 s 0 33819 28 33867 4 wl1_84
port 105 nsew
rlabel metal2 s 0 34293 28 34341 4 wl0_85
port 106 nsew
rlabel metal2 s 0 34073 28 34121 4 wl1_85
port 107 nsew
rlabel metal2 s 0 34389 28 34437 4 wl0_86
port 108 nsew
rlabel metal2 s 0 34609 28 34657 4 wl1_86
port 109 nsew
rlabel metal2 s 0 35083 28 35131 4 wl0_87
port 110 nsew
rlabel metal2 s 0 34863 28 34911 4 wl1_87
port 111 nsew
rlabel metal2 s 0 35179 28 35227 4 wl0_88
port 112 nsew
rlabel metal2 s 0 35399 28 35447 4 wl1_88
port 113 nsew
rlabel metal2 s 0 35873 28 35921 4 wl0_89
port 114 nsew
rlabel metal2 s 0 35653 28 35701 4 wl1_89
port 115 nsew
rlabel metal2 s 0 35969 28 36017 4 wl0_90
port 116 nsew
rlabel metal2 s 0 36189 28 36237 4 wl1_90
port 117 nsew
rlabel metal2 s 0 36663 28 36711 4 wl0_91
port 118 nsew
rlabel metal2 s 0 36443 28 36491 4 wl1_91
port 119 nsew
rlabel metal2 s 0 36759 28 36807 4 wl0_92
port 120 nsew
rlabel metal2 s 0 36979 28 37027 4 wl1_92
port 121 nsew
rlabel metal2 s 0 37453 28 37501 4 wl0_93
port 122 nsew
rlabel metal2 s 0 37233 28 37281 4 wl1_93
port 123 nsew
rlabel metal2 s 0 37549 28 37597 4 wl0_94
port 124 nsew
rlabel metal2 s 0 37769 28 37817 4 wl1_94
port 125 nsew
rlabel metal2 s 0 38243 28 38291 4 wl0_95
port 126 nsew
rlabel metal2 s 0 38023 28 38071 4 wl1_95
port 127 nsew
rlabel metal2 s 0 38339 28 38387 4 wl0_96
port 128 nsew
rlabel metal2 s 0 38559 28 38607 4 wl1_96
port 129 nsew
rlabel metal2 s 0 13753 28 13801 4 wl0_33
port 130 nsew
rlabel metal2 s 0 13533 28 13581 4 wl1_33
port 131 nsew
rlabel metal2 s 0 13849 28 13897 4 wl0_34
port 132 nsew
rlabel metal2 s 0 14069 28 14117 4 wl1_34
port 133 nsew
rlabel metal2 s 0 14543 28 14591 4 wl0_35
port 134 nsew
rlabel metal2 s 0 14323 28 14371 4 wl1_35
port 135 nsew
rlabel metal2 s 0 14639 28 14687 4 wl0_36
port 136 nsew
rlabel metal2 s 0 14859 28 14907 4 wl1_36
port 137 nsew
rlabel metal2 s 0 15333 28 15381 4 wl0_37
port 138 nsew
rlabel metal2 s 0 15113 28 15161 4 wl1_37
port 139 nsew
rlabel metal2 s 0 15429 28 15477 4 wl0_38
port 140 nsew
rlabel metal2 s 0 15649 28 15697 4 wl1_38
port 141 nsew
rlabel metal2 s 0 16123 28 16171 4 wl0_39
port 142 nsew
rlabel metal2 s 0 15903 28 15951 4 wl1_39
port 143 nsew
rlabel metal2 s 0 16219 28 16267 4 wl0_40
port 144 nsew
rlabel metal2 s 0 16439 28 16487 4 wl1_40
port 145 nsew
rlabel metal2 s 0 16913 28 16961 4 wl0_41
port 146 nsew
rlabel metal2 s 0 16693 28 16741 4 wl1_41
port 147 nsew
rlabel metal2 s 0 17009 28 17057 4 wl0_42
port 148 nsew
rlabel metal2 s 0 17229 28 17277 4 wl1_42
port 149 nsew
rlabel metal2 s 0 17703 28 17751 4 wl0_43
port 150 nsew
rlabel metal2 s 0 17483 28 17531 4 wl1_43
port 151 nsew
rlabel metal2 s 0 17799 28 17847 4 wl0_44
port 152 nsew
rlabel metal2 s 0 18019 28 18067 4 wl1_44
port 153 nsew
rlabel metal2 s 0 18493 28 18541 4 wl0_45
port 154 nsew
rlabel metal2 s 0 18273 28 18321 4 wl1_45
port 155 nsew
rlabel metal2 s 0 18589 28 18637 4 wl0_46
port 156 nsew
rlabel metal2 s 0 18809 28 18857 4 wl1_46
port 157 nsew
rlabel metal2 s 0 19283 28 19331 4 wl0_47
port 158 nsew
rlabel metal2 s 0 19063 28 19111 4 wl1_47
port 159 nsew
rlabel metal2 s 0 19379 28 19427 4 wl0_48
port 160 nsew
rlabel metal2 s 0 19599 28 19647 4 wl1_48
port 161 nsew
rlabel metal2 s 0 20073 28 20121 4 wl0_49
port 162 nsew
rlabel metal2 s 0 19853 28 19901 4 wl1_49
port 163 nsew
rlabel metal2 s 0 20169 28 20217 4 wl0_50
port 164 nsew
rlabel metal2 s 0 20389 28 20437 4 wl1_50
port 165 nsew
rlabel metal2 s 0 20863 28 20911 4 wl0_51
port 166 nsew
rlabel metal2 s 0 20643 28 20691 4 wl1_51
port 167 nsew
rlabel metal2 s 0 20959 28 21007 4 wl0_52
port 168 nsew
rlabel metal2 s 0 21179 28 21227 4 wl1_52
port 169 nsew
rlabel metal2 s 0 21653 28 21701 4 wl0_53
port 170 nsew
rlabel metal2 s 0 21433 28 21481 4 wl1_53
port 171 nsew
rlabel metal2 s 0 21749 28 21797 4 wl0_54
port 172 nsew
rlabel metal2 s 0 21969 28 22017 4 wl1_54
port 173 nsew
rlabel metal2 s 0 22443 28 22491 4 wl0_55
port 174 nsew
rlabel metal2 s 0 22223 28 22271 4 wl1_55
port 175 nsew
rlabel metal2 s 0 22539 28 22587 4 wl0_56
port 176 nsew
rlabel metal2 s 0 22759 28 22807 4 wl1_56
port 177 nsew
rlabel metal2 s 0 23233 28 23281 4 wl0_57
port 178 nsew
rlabel metal2 s 0 23013 28 23061 4 wl1_57
port 179 nsew
rlabel metal2 s 0 23329 28 23377 4 wl0_58
port 180 nsew
rlabel metal2 s 0 23549 28 23597 4 wl1_58
port 181 nsew
rlabel metal2 s 0 24023 28 24071 4 wl0_59
port 182 nsew
rlabel metal2 s 0 23803 28 23851 4 wl1_59
port 183 nsew
rlabel metal2 s 0 24119 28 24167 4 wl0_60
port 184 nsew
rlabel metal2 s 0 24339 28 24387 4 wl1_60
port 185 nsew
rlabel metal2 s 0 24813 28 24861 4 wl0_61
port 186 nsew
rlabel metal2 s 0 24593 28 24641 4 wl1_61
port 187 nsew
rlabel metal2 s 0 24909 28 24957 4 wl0_62
port 188 nsew
rlabel metal2 s 0 25129 28 25177 4 wl1_62
port 189 nsew
rlabel metal2 s 0 25603 28 25651 4 wl0_63
port 190 nsew
rlabel metal2 s 0 25383 28 25431 4 wl1_63
port 191 nsew
rlabel metal2 s 0 25699 28 25747 4 wl0_64
port 192 nsew
rlabel metal2 s 0 25919 28 25967 4 wl1_64
port 193 nsew
rlabel metal2 s 0 1113 28 1161 4 wl0_1
port 194 nsew
rlabel metal2 s 0 893 28 941 4 wl1_1
port 195 nsew
rlabel metal2 s 0 1209 28 1257 4 wl0_2
port 196 nsew
rlabel metal2 s 0 1429 28 1477 4 wl1_2
port 197 nsew
rlabel metal2 s 0 1903 28 1951 4 wl0_3
port 198 nsew
rlabel metal2 s 0 1683 28 1731 4 wl1_3
port 199 nsew
rlabel metal2 s 0 1999 28 2047 4 wl0_4
port 200 nsew
rlabel metal2 s 0 2219 28 2267 4 wl1_4
port 201 nsew
rlabel metal2 s 0 2693 28 2741 4 wl0_5
port 202 nsew
rlabel metal2 s 0 2473 28 2521 4 wl1_5
port 203 nsew
rlabel metal2 s 0 2789 28 2837 4 wl0_6
port 204 nsew
rlabel metal2 s 0 3009 28 3057 4 wl1_6
port 205 nsew
rlabel metal2 s 0 3483 28 3531 4 wl0_7
port 206 nsew
rlabel metal2 s 0 3263 28 3311 4 wl1_7
port 207 nsew
rlabel metal2 s 0 3579 28 3627 4 wl0_8
port 208 nsew
rlabel metal2 s 0 3799 28 3847 4 wl1_8
port 209 nsew
rlabel metal2 s 0 4273 28 4321 4 wl0_9
port 210 nsew
rlabel metal2 s 0 4053 28 4101 4 wl1_9
port 211 nsew
rlabel metal2 s 0 4369 28 4417 4 wl0_10
port 212 nsew
rlabel metal2 s 0 4589 28 4637 4 wl1_10
port 213 nsew
rlabel metal2 s 0 5063 28 5111 4 wl0_11
port 214 nsew
rlabel metal2 s 0 4843 28 4891 4 wl1_11
port 215 nsew
rlabel metal2 s 0 5159 28 5207 4 wl0_12
port 216 nsew
rlabel metal2 s 0 5379 28 5427 4 wl1_12
port 217 nsew
rlabel metal2 s 0 5853 28 5901 4 wl0_13
port 218 nsew
rlabel metal2 s 0 5633 28 5681 4 wl1_13
port 219 nsew
rlabel metal2 s 0 5949 28 5997 4 wl0_14
port 220 nsew
rlabel metal2 s 0 6169 28 6217 4 wl1_14
port 221 nsew
rlabel metal2 s 0 6643 28 6691 4 wl0_15
port 222 nsew
rlabel metal2 s 0 6423 28 6471 4 wl1_15
port 223 nsew
rlabel metal2 s 0 6739 28 6787 4 wl0_16
port 224 nsew
rlabel metal2 s 0 6959 28 7007 4 wl1_16
port 225 nsew
rlabel metal2 s 0 7433 28 7481 4 wl0_17
port 226 nsew
rlabel metal2 s 0 7213 28 7261 4 wl1_17
port 227 nsew
rlabel metal2 s 0 7529 28 7577 4 wl0_18
port 228 nsew
rlabel metal2 s 0 7749 28 7797 4 wl1_18
port 229 nsew
rlabel metal2 s 0 8223 28 8271 4 wl0_19
port 230 nsew
rlabel metal2 s 0 8003 28 8051 4 wl1_19
port 231 nsew
rlabel metal2 s 0 8319 28 8367 4 wl0_20
port 232 nsew
rlabel metal2 s 0 8539 28 8587 4 wl1_20
port 233 nsew
rlabel metal2 s 0 9013 28 9061 4 wl0_21
port 234 nsew
rlabel metal2 s 0 8793 28 8841 4 wl1_21
port 235 nsew
rlabel metal2 s 0 9109 28 9157 4 wl0_22
port 236 nsew
rlabel metal2 s 0 9329 28 9377 4 wl1_22
port 237 nsew
rlabel metal2 s 0 9803 28 9851 4 wl0_23
port 238 nsew
rlabel metal2 s 0 9583 28 9631 4 wl1_23
port 239 nsew
rlabel metal2 s 0 9899 28 9947 4 wl0_24
port 240 nsew
rlabel metal2 s 0 10119 28 10167 4 wl1_24
port 241 nsew
rlabel metal2 s 0 10593 28 10641 4 wl0_25
port 242 nsew
rlabel metal2 s 0 10373 28 10421 4 wl1_25
port 243 nsew
rlabel metal2 s 0 10689 28 10737 4 wl0_26
port 244 nsew
rlabel metal2 s 0 10909 28 10957 4 wl1_26
port 245 nsew
rlabel metal2 s 0 11383 28 11431 4 wl0_27
port 246 nsew
rlabel metal2 s 0 11163 28 11211 4 wl1_27
port 247 nsew
rlabel metal2 s 0 11479 28 11527 4 wl0_28
port 248 nsew
rlabel metal2 s 0 11699 28 11747 4 wl1_28
port 249 nsew
rlabel metal2 s 0 12173 28 12221 4 wl0_29
port 250 nsew
rlabel metal2 s 0 11953 28 12001 4 wl1_29
port 251 nsew
rlabel metal2 s 0 12269 28 12317 4 wl0_30
port 252 nsew
rlabel metal2 s 0 12489 28 12537 4 wl1_30
port 253 nsew
rlabel metal2 s 0 12963 28 13011 4 wl0_31
port 254 nsew
rlabel metal2 s 0 12743 28 12791 4 wl1_31
port 255 nsew
rlabel metal2 s 0 13059 28 13107 4 wl0_32
port 256 nsew
rlabel metal2 s 0 13279 28 13327 4 wl1_32
port 257 nsew
<< properties >>
string FIXED_BBOX 0 0 624 51745
string GDS_END 1246178
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 1137428
<< end >>

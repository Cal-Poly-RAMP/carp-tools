magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< poly >>
rect 1671 435 1701 1392
rect 2295 559 2325 1392
rect 2919 683 2949 1392
rect 3543 807 3573 1392
rect 4167 931 4197 1392
rect 4791 1055 4821 1392
rect 5415 1179 5445 1392
rect 6039 1303 6069 1392
rect 6021 1287 6087 1303
rect 6021 1253 6037 1287
rect 6071 1253 6087 1287
rect 6021 1237 6087 1253
rect 5397 1163 5463 1179
rect 5397 1129 5413 1163
rect 5447 1129 5463 1163
rect 5397 1113 5463 1129
rect 4773 1039 4839 1055
rect 4773 1005 4789 1039
rect 4823 1005 4839 1039
rect 4773 989 4839 1005
rect 4149 915 4215 931
rect 4149 881 4165 915
rect 4199 881 4215 915
rect 4149 865 4215 881
rect 3525 791 3591 807
rect 3525 757 3541 791
rect 3575 757 3591 791
rect 3525 741 3591 757
rect 2901 667 2967 683
rect 2901 633 2917 667
rect 2951 633 2967 667
rect 2901 617 2967 633
rect 2277 543 2343 559
rect 2277 509 2293 543
rect 2327 509 2343 543
rect 2277 493 2343 509
rect 6663 435 6693 1392
rect 7287 559 7317 1392
rect 7911 683 7941 1392
rect 8535 807 8565 1392
rect 9159 931 9189 1392
rect 9783 1055 9813 1392
rect 10407 1179 10437 1392
rect 11031 1303 11061 1392
rect 11013 1287 11079 1303
rect 11013 1253 11029 1287
rect 11063 1253 11079 1287
rect 11013 1237 11079 1253
rect 10389 1163 10455 1179
rect 10389 1129 10405 1163
rect 10439 1129 10455 1163
rect 10389 1113 10455 1129
rect 9765 1039 9831 1055
rect 9765 1005 9781 1039
rect 9815 1005 9831 1039
rect 9765 989 9831 1005
rect 9141 915 9207 931
rect 9141 881 9157 915
rect 9191 881 9207 915
rect 9141 865 9207 881
rect 8517 791 8583 807
rect 8517 757 8533 791
rect 8567 757 8583 791
rect 8517 741 8583 757
rect 7893 667 7959 683
rect 7893 633 7909 667
rect 7943 633 7959 667
rect 7893 617 7959 633
rect 7269 543 7335 559
rect 7269 509 7285 543
rect 7319 509 7335 543
rect 7269 493 7335 509
rect 11655 435 11685 1392
rect 12279 559 12309 1392
rect 12903 683 12933 1392
rect 13527 807 13557 1392
rect 14151 931 14181 1392
rect 14775 1055 14805 1392
rect 15399 1179 15429 1392
rect 16023 1303 16053 1392
rect 16005 1287 16071 1303
rect 16005 1253 16021 1287
rect 16055 1253 16071 1287
rect 16005 1237 16071 1253
rect 15381 1163 15447 1179
rect 15381 1129 15397 1163
rect 15431 1129 15447 1163
rect 15381 1113 15447 1129
rect 14757 1039 14823 1055
rect 14757 1005 14773 1039
rect 14807 1005 14823 1039
rect 14757 989 14823 1005
rect 14133 915 14199 931
rect 14133 881 14149 915
rect 14183 881 14199 915
rect 14133 865 14199 881
rect 13509 791 13575 807
rect 13509 757 13525 791
rect 13559 757 13575 791
rect 13509 741 13575 757
rect 12885 667 12951 683
rect 12885 633 12901 667
rect 12935 633 12951 667
rect 12885 617 12951 633
rect 12261 543 12327 559
rect 12261 509 12277 543
rect 12311 509 12327 543
rect 12261 493 12327 509
rect 16647 435 16677 1392
rect 17271 559 17301 1392
rect 17895 683 17925 1392
rect 18519 807 18549 1392
rect 19143 931 19173 1392
rect 19767 1055 19797 1392
rect 20391 1179 20421 1392
rect 21015 1303 21045 1392
rect 20997 1287 21063 1303
rect 20997 1253 21013 1287
rect 21047 1253 21063 1287
rect 20997 1237 21063 1253
rect 20373 1163 20439 1179
rect 20373 1129 20389 1163
rect 20423 1129 20439 1163
rect 20373 1113 20439 1129
rect 19749 1039 19815 1055
rect 19749 1005 19765 1039
rect 19799 1005 19815 1039
rect 19749 989 19815 1005
rect 19125 915 19191 931
rect 19125 881 19141 915
rect 19175 881 19191 915
rect 19125 865 19191 881
rect 18501 791 18567 807
rect 18501 757 18517 791
rect 18551 757 18567 791
rect 18501 741 18567 757
rect 17877 667 17943 683
rect 17877 633 17893 667
rect 17927 633 17943 667
rect 17877 617 17943 633
rect 17253 543 17319 559
rect 17253 509 17269 543
rect 17303 509 17319 543
rect 17253 493 17319 509
rect 21639 435 21669 1392
rect 22263 559 22293 1392
rect 22887 683 22917 1392
rect 23511 807 23541 1392
rect 24135 931 24165 1392
rect 24759 1055 24789 1392
rect 25383 1179 25413 1392
rect 26007 1303 26037 1392
rect 25989 1287 26055 1303
rect 25989 1253 26005 1287
rect 26039 1253 26055 1287
rect 25989 1237 26055 1253
rect 25365 1163 25431 1179
rect 25365 1129 25381 1163
rect 25415 1129 25431 1163
rect 25365 1113 25431 1129
rect 24741 1039 24807 1055
rect 24741 1005 24757 1039
rect 24791 1005 24807 1039
rect 24741 989 24807 1005
rect 24117 915 24183 931
rect 24117 881 24133 915
rect 24167 881 24183 915
rect 24117 865 24183 881
rect 23493 791 23559 807
rect 23493 757 23509 791
rect 23543 757 23559 791
rect 23493 741 23559 757
rect 22869 667 22935 683
rect 22869 633 22885 667
rect 22919 633 22935 667
rect 22869 617 22935 633
rect 22245 543 22311 559
rect 22245 509 22261 543
rect 22295 509 22311 543
rect 22245 493 22311 509
rect 26631 435 26661 1392
rect 27255 559 27285 1392
rect 27879 683 27909 1392
rect 28503 807 28533 1392
rect 29127 931 29157 1392
rect 29751 1055 29781 1392
rect 30375 1179 30405 1392
rect 30999 1303 31029 1392
rect 30981 1287 31047 1303
rect 30981 1253 30997 1287
rect 31031 1253 31047 1287
rect 30981 1237 31047 1253
rect 30357 1163 30423 1179
rect 30357 1129 30373 1163
rect 30407 1129 30423 1163
rect 30357 1113 30423 1129
rect 29733 1039 29799 1055
rect 29733 1005 29749 1039
rect 29783 1005 29799 1039
rect 29733 989 29799 1005
rect 29109 915 29175 931
rect 29109 881 29125 915
rect 29159 881 29175 915
rect 29109 865 29175 881
rect 28485 791 28551 807
rect 28485 757 28501 791
rect 28535 757 28551 791
rect 28485 741 28551 757
rect 27861 667 27927 683
rect 27861 633 27877 667
rect 27911 633 27927 667
rect 27861 617 27927 633
rect 27237 543 27303 559
rect 27237 509 27253 543
rect 27287 509 27303 543
rect 27237 493 27303 509
rect 31623 435 31653 1392
rect 32247 559 32277 1392
rect 32871 683 32901 1392
rect 33495 807 33525 1392
rect 34119 931 34149 1392
rect 34743 1055 34773 1392
rect 35367 1179 35397 1392
rect 35991 1303 36021 1392
rect 35973 1287 36039 1303
rect 35973 1253 35989 1287
rect 36023 1253 36039 1287
rect 35973 1237 36039 1253
rect 35349 1163 35415 1179
rect 35349 1129 35365 1163
rect 35399 1129 35415 1163
rect 35349 1113 35415 1129
rect 34725 1039 34791 1055
rect 34725 1005 34741 1039
rect 34775 1005 34791 1039
rect 34725 989 34791 1005
rect 34101 915 34167 931
rect 34101 881 34117 915
rect 34151 881 34167 915
rect 34101 865 34167 881
rect 33477 791 33543 807
rect 33477 757 33493 791
rect 33527 757 33543 791
rect 33477 741 33543 757
rect 32853 667 32919 683
rect 32853 633 32869 667
rect 32903 633 32919 667
rect 32853 617 32919 633
rect 32229 543 32295 559
rect 32229 509 32245 543
rect 32279 509 32295 543
rect 32229 493 32295 509
rect 36615 435 36645 1392
rect 37239 559 37269 1392
rect 37863 683 37893 1392
rect 38487 807 38517 1392
rect 39111 931 39141 1392
rect 39735 1055 39765 1392
rect 40359 1179 40389 1392
rect 40983 1303 41013 1392
rect 40965 1287 41031 1303
rect 40965 1253 40981 1287
rect 41015 1253 41031 1287
rect 40965 1237 41031 1253
rect 40341 1163 40407 1179
rect 40341 1129 40357 1163
rect 40391 1129 40407 1163
rect 40341 1113 40407 1129
rect 39717 1039 39783 1055
rect 39717 1005 39733 1039
rect 39767 1005 39783 1039
rect 39717 989 39783 1005
rect 39093 915 39159 931
rect 39093 881 39109 915
rect 39143 881 39159 915
rect 39093 865 39159 881
rect 38469 791 38535 807
rect 38469 757 38485 791
rect 38519 757 38535 791
rect 38469 741 38535 757
rect 37845 667 37911 683
rect 37845 633 37861 667
rect 37895 633 37911 667
rect 37845 617 37911 633
rect 37221 543 37287 559
rect 37221 509 37237 543
rect 37271 509 37287 543
rect 37221 493 37287 509
rect 1653 419 1719 435
rect 1653 385 1669 419
rect 1703 385 1719 419
rect 1653 369 1719 385
rect 6645 419 6711 435
rect 6645 385 6661 419
rect 6695 385 6711 419
rect 6645 369 6711 385
rect 11637 419 11703 435
rect 11637 385 11653 419
rect 11687 385 11703 419
rect 11637 369 11703 385
rect 16629 419 16695 435
rect 16629 385 16645 419
rect 16679 385 16695 419
rect 16629 369 16695 385
rect 21621 419 21687 435
rect 21621 385 21637 419
rect 21671 385 21687 419
rect 21621 369 21687 385
rect 26613 419 26679 435
rect 26613 385 26629 419
rect 26663 385 26679 419
rect 26613 369 26679 385
rect 31605 419 31671 435
rect 31605 385 31621 419
rect 31655 385 31671 419
rect 31605 369 31671 385
rect 36597 419 36663 435
rect 36597 385 36613 419
rect 36647 385 36663 419
rect 36597 369 36663 385
<< polycont >>
rect 6037 1253 6071 1287
rect 5413 1129 5447 1163
rect 4789 1005 4823 1039
rect 4165 881 4199 915
rect 3541 757 3575 791
rect 2917 633 2951 667
rect 2293 509 2327 543
rect 11029 1253 11063 1287
rect 10405 1129 10439 1163
rect 9781 1005 9815 1039
rect 9157 881 9191 915
rect 8533 757 8567 791
rect 7909 633 7943 667
rect 7285 509 7319 543
rect 16021 1253 16055 1287
rect 15397 1129 15431 1163
rect 14773 1005 14807 1039
rect 14149 881 14183 915
rect 13525 757 13559 791
rect 12901 633 12935 667
rect 12277 509 12311 543
rect 21013 1253 21047 1287
rect 20389 1129 20423 1163
rect 19765 1005 19799 1039
rect 19141 881 19175 915
rect 18517 757 18551 791
rect 17893 633 17927 667
rect 17269 509 17303 543
rect 26005 1253 26039 1287
rect 25381 1129 25415 1163
rect 24757 1005 24791 1039
rect 24133 881 24167 915
rect 23509 757 23543 791
rect 22885 633 22919 667
rect 22261 509 22295 543
rect 30997 1253 31031 1287
rect 30373 1129 30407 1163
rect 29749 1005 29783 1039
rect 29125 881 29159 915
rect 28501 757 28535 791
rect 27877 633 27911 667
rect 27253 509 27287 543
rect 35989 1253 36023 1287
rect 35365 1129 35399 1163
rect 34741 1005 34775 1039
rect 34117 881 34151 915
rect 33493 757 33527 791
rect 32869 633 32903 667
rect 32245 509 32279 543
rect 40981 1253 41015 1287
rect 40357 1129 40391 1163
rect 39733 1005 39767 1039
rect 39109 881 39143 915
rect 38485 757 38519 791
rect 37861 633 37895 667
rect 37237 509 37271 543
rect 1669 385 1703 419
rect 6661 385 6695 419
rect 11653 385 11687 419
rect 16645 385 16679 419
rect 21637 385 21671 419
rect 26629 385 26663 419
rect 31621 385 31655 419
rect 36613 385 36647 419
<< locali >>
rect 6037 1287 6071 1303
rect 6037 1237 6071 1253
rect 11029 1287 11063 1303
rect 11029 1237 11063 1253
rect 16021 1287 16055 1303
rect 16021 1237 16055 1253
rect 21013 1287 21047 1303
rect 21013 1237 21047 1253
rect 26005 1287 26039 1303
rect 26005 1237 26039 1253
rect 30997 1287 31031 1303
rect 30997 1237 31031 1253
rect 35989 1287 36023 1303
rect 35989 1237 36023 1253
rect 40981 1287 41015 1303
rect 40981 1237 41015 1253
rect 5413 1163 5447 1179
rect 5413 1113 5447 1129
rect 10405 1163 10439 1179
rect 10405 1113 10439 1129
rect 15397 1163 15431 1179
rect 15397 1113 15431 1129
rect 20389 1163 20423 1179
rect 20389 1113 20423 1129
rect 25381 1163 25415 1179
rect 25381 1113 25415 1129
rect 30373 1163 30407 1179
rect 30373 1113 30407 1129
rect 35365 1163 35399 1179
rect 35365 1113 35399 1129
rect 40357 1163 40391 1179
rect 40357 1113 40391 1129
rect 4789 1039 4823 1055
rect 4789 989 4823 1005
rect 9781 1039 9815 1055
rect 9781 989 9815 1005
rect 14773 1039 14807 1055
rect 14773 989 14807 1005
rect 19765 1039 19799 1055
rect 19765 989 19799 1005
rect 24757 1039 24791 1055
rect 24757 989 24791 1005
rect 29749 1039 29783 1055
rect 29749 989 29783 1005
rect 34741 1039 34775 1055
rect 34741 989 34775 1005
rect 39733 1039 39767 1055
rect 39733 989 39767 1005
rect 4165 915 4199 931
rect 4165 865 4199 881
rect 9157 915 9191 931
rect 9157 865 9191 881
rect 14149 915 14183 931
rect 14149 865 14183 881
rect 19141 915 19175 931
rect 19141 865 19175 881
rect 24133 915 24167 931
rect 24133 865 24167 881
rect 29125 915 29159 931
rect 29125 865 29159 881
rect 34117 915 34151 931
rect 34117 865 34151 881
rect 39109 915 39143 931
rect 39109 865 39143 881
rect 3541 791 3575 807
rect 3541 741 3575 757
rect 8533 791 8567 807
rect 8533 741 8567 757
rect 13525 791 13559 807
rect 13525 741 13559 757
rect 18517 791 18551 807
rect 18517 741 18551 757
rect 23509 791 23543 807
rect 23509 741 23543 757
rect 28501 791 28535 807
rect 28501 741 28535 757
rect 33493 791 33527 807
rect 33493 741 33527 757
rect 38485 791 38519 807
rect 38485 741 38519 757
rect 2917 667 2951 683
rect 2917 617 2951 633
rect 7909 667 7943 683
rect 7909 617 7943 633
rect 12901 667 12935 683
rect 12901 617 12935 633
rect 17893 667 17927 683
rect 17893 617 17927 633
rect 22885 667 22919 683
rect 22885 617 22919 633
rect 27877 667 27911 683
rect 27877 617 27911 633
rect 32869 667 32903 683
rect 32869 617 32903 633
rect 37861 667 37895 683
rect 37861 617 37895 633
rect 2293 543 2327 559
rect 2293 493 2327 509
rect 7285 543 7319 559
rect 7285 493 7319 509
rect 12277 543 12311 559
rect 12277 493 12311 509
rect 17269 543 17303 559
rect 17269 493 17303 509
rect 22261 543 22295 559
rect 22261 493 22295 509
rect 27253 543 27287 559
rect 27253 493 27287 509
rect 32245 543 32279 559
rect 32245 493 32279 509
rect 37237 543 37271 559
rect 37237 493 37271 509
rect 1669 419 1703 435
rect 1669 369 1703 385
rect 6661 419 6695 435
rect 6661 369 6695 385
rect 11653 419 11687 435
rect 11653 369 11687 385
rect 16645 419 16679 435
rect 16645 369 16679 385
rect 21637 419 21671 435
rect 21637 369 21671 385
rect 26629 419 26663 435
rect 26629 369 26663 385
rect 31621 419 31655 435
rect 31621 369 31655 385
rect 36613 419 36647 435
rect 36613 369 36647 385
<< viali >>
rect 6037 1253 6071 1287
rect 11029 1253 11063 1287
rect 16021 1253 16055 1287
rect 21013 1253 21047 1287
rect 26005 1253 26039 1287
rect 30997 1253 31031 1287
rect 35989 1253 36023 1287
rect 40981 1253 41015 1287
rect 5413 1129 5447 1163
rect 10405 1129 10439 1163
rect 15397 1129 15431 1163
rect 20389 1129 20423 1163
rect 25381 1129 25415 1163
rect 30373 1129 30407 1163
rect 35365 1129 35399 1163
rect 40357 1129 40391 1163
rect 4789 1005 4823 1039
rect 9781 1005 9815 1039
rect 14773 1005 14807 1039
rect 19765 1005 19799 1039
rect 24757 1005 24791 1039
rect 29749 1005 29783 1039
rect 34741 1005 34775 1039
rect 39733 1005 39767 1039
rect 4165 881 4199 915
rect 9157 881 9191 915
rect 14149 881 14183 915
rect 19141 881 19175 915
rect 24133 881 24167 915
rect 29125 881 29159 915
rect 34117 881 34151 915
rect 39109 881 39143 915
rect 3541 757 3575 791
rect 8533 757 8567 791
rect 13525 757 13559 791
rect 18517 757 18551 791
rect 23509 757 23543 791
rect 28501 757 28535 791
rect 33493 757 33527 791
rect 38485 757 38519 791
rect 2917 633 2951 667
rect 7909 633 7943 667
rect 12901 633 12935 667
rect 17893 633 17927 667
rect 22885 633 22919 667
rect 27877 633 27911 667
rect 32869 633 32903 667
rect 37861 633 37895 667
rect 2293 509 2327 543
rect 7285 509 7319 543
rect 12277 509 12311 543
rect 17269 509 17303 543
rect 22261 509 22295 543
rect 27253 509 27287 543
rect 32245 509 32279 543
rect 37237 509 37271 543
rect 1669 385 1703 419
rect 6661 385 6695 419
rect 11653 385 11687 419
rect 16645 385 16679 419
rect 21637 385 21671 419
rect 26629 385 26663 419
rect 31621 385 31655 419
rect 36613 385 36647 419
<< metal1 >>
rect 1454 2624 1482 2680
rect 1918 2624 1946 2680
rect 2050 2624 2078 2680
rect 2514 2624 2542 2680
rect 2702 2624 2730 2680
rect 3166 2624 3194 2680
rect 3298 2624 3326 2680
rect 3762 2624 3790 2680
rect 3950 2624 3978 2680
rect 4414 2624 4442 2680
rect 4546 2624 4574 2680
rect 5010 2624 5038 2680
rect 5198 2624 5226 2680
rect 5662 2624 5690 2680
rect 5794 2624 5822 2680
rect 6258 2624 6286 2680
rect 6446 2624 6474 2680
rect 6910 2624 6938 2680
rect 7042 2624 7070 2680
rect 7506 2624 7534 2680
rect 7694 2624 7722 2680
rect 8158 2624 8186 2680
rect 8290 2624 8318 2680
rect 8754 2624 8782 2680
rect 8942 2624 8970 2680
rect 9406 2624 9434 2680
rect 9538 2624 9566 2680
rect 10002 2624 10030 2680
rect 10190 2624 10218 2680
rect 10654 2624 10682 2680
rect 10786 2624 10814 2680
rect 11250 2624 11278 2680
rect 11438 2624 11466 2680
rect 11902 2624 11930 2680
rect 12034 2624 12062 2680
rect 12498 2624 12526 2680
rect 12686 2624 12714 2680
rect 13150 2624 13178 2680
rect 13282 2624 13310 2680
rect 13746 2624 13774 2680
rect 13934 2624 13962 2680
rect 14398 2624 14426 2680
rect 14530 2624 14558 2680
rect 14994 2624 15022 2680
rect 15182 2624 15210 2680
rect 15646 2624 15674 2680
rect 15778 2624 15806 2680
rect 16242 2624 16270 2680
rect 16430 2624 16458 2680
rect 16894 2624 16922 2680
rect 17026 2624 17054 2680
rect 17490 2624 17518 2680
rect 17678 2624 17706 2680
rect 18142 2624 18170 2680
rect 18274 2624 18302 2680
rect 18738 2624 18766 2680
rect 18926 2624 18954 2680
rect 19390 2624 19418 2680
rect 19522 2624 19550 2680
rect 19986 2624 20014 2680
rect 20174 2624 20202 2680
rect 20638 2624 20666 2680
rect 20770 2624 20798 2680
rect 21234 2624 21262 2680
rect 21422 2624 21450 2680
rect 21886 2624 21914 2680
rect 22018 2624 22046 2680
rect 22482 2624 22510 2680
rect 22670 2624 22698 2680
rect 23134 2624 23162 2680
rect 23266 2624 23294 2680
rect 23730 2624 23758 2680
rect 23918 2624 23946 2680
rect 24382 2624 24410 2680
rect 24514 2624 24542 2680
rect 24978 2624 25006 2680
rect 25166 2624 25194 2680
rect 25630 2624 25658 2680
rect 25762 2624 25790 2680
rect 26226 2624 26254 2680
rect 26414 2624 26442 2680
rect 26878 2624 26906 2680
rect 27010 2624 27038 2680
rect 27474 2624 27502 2680
rect 27662 2624 27690 2680
rect 28126 2624 28154 2680
rect 28258 2624 28286 2680
rect 28722 2624 28750 2680
rect 28910 2624 28938 2680
rect 29374 2624 29402 2680
rect 29506 2624 29534 2680
rect 29970 2624 29998 2680
rect 30158 2624 30186 2680
rect 30622 2624 30650 2680
rect 30754 2624 30782 2680
rect 31218 2624 31246 2680
rect 31406 2624 31434 2680
rect 31870 2624 31898 2680
rect 32002 2624 32030 2680
rect 32466 2624 32494 2680
rect 32654 2624 32682 2680
rect 33118 2624 33146 2680
rect 33250 2624 33278 2680
rect 33714 2624 33742 2680
rect 33902 2624 33930 2680
rect 34366 2624 34394 2680
rect 34498 2624 34526 2680
rect 34962 2624 34990 2680
rect 35150 2624 35178 2680
rect 35614 2624 35642 2680
rect 35746 2624 35774 2680
rect 36210 2624 36238 2680
rect 36398 2624 36426 2680
rect 36862 2624 36890 2680
rect 36994 2624 37022 2680
rect 37458 2624 37486 2680
rect 37646 2624 37674 2680
rect 38110 2624 38138 2680
rect 38242 2624 38270 2680
rect 38706 2624 38734 2680
rect 38894 2624 38922 2680
rect 39358 2624 39386 2680
rect 39490 2624 39518 2680
rect 39954 2624 39982 2680
rect 40142 2624 40170 2680
rect 40606 2624 40634 2680
rect 40738 2624 40766 2680
rect 41202 2624 41230 2680
rect 1454 274 1482 1364
rect 1654 376 1660 428
rect 1712 376 1718 428
rect 1436 222 1442 274
rect 1494 222 1500 274
rect 1918 150 1946 1364
rect 2050 150 2078 1364
rect 2278 500 2284 552
rect 2336 500 2342 552
rect 2514 274 2542 1364
rect 2702 274 2730 1364
rect 2902 624 2908 676
rect 2960 624 2966 676
rect 2496 222 2502 274
rect 2554 222 2560 274
rect 2684 222 2690 274
rect 2742 222 2748 274
rect 3166 150 3194 1364
rect 3298 150 3326 1364
rect 3526 748 3532 800
rect 3584 748 3590 800
rect 3762 274 3790 1364
rect 3950 274 3978 1364
rect 4150 872 4156 924
rect 4208 872 4214 924
rect 3744 222 3750 274
rect 3802 222 3808 274
rect 3932 222 3938 274
rect 3990 222 3996 274
rect 4414 150 4442 1364
rect 4546 150 4574 1364
rect 4774 996 4780 1048
rect 4832 996 4838 1048
rect 5010 274 5038 1364
rect 5198 274 5226 1364
rect 5398 1120 5404 1172
rect 5456 1120 5462 1172
rect 4992 222 4998 274
rect 5050 222 5056 274
rect 5180 222 5186 274
rect 5238 222 5244 274
rect 5662 150 5690 1364
rect 5794 150 5822 1364
rect 6022 1244 6028 1296
rect 6080 1244 6086 1296
rect 6258 274 6286 1364
rect 6446 274 6474 1364
rect 6646 376 6652 428
rect 6704 376 6710 428
rect 6240 222 6246 274
rect 6298 222 6304 274
rect 6428 222 6434 274
rect 6486 222 6492 274
rect 6910 150 6938 1364
rect 7042 150 7070 1364
rect 7270 500 7276 552
rect 7328 500 7334 552
rect 7506 274 7534 1364
rect 7694 274 7722 1364
rect 7894 624 7900 676
rect 7952 624 7958 676
rect 7488 222 7494 274
rect 7546 222 7552 274
rect 7676 222 7682 274
rect 7734 222 7740 274
rect 8158 150 8186 1364
rect 8290 150 8318 1364
rect 8518 748 8524 800
rect 8576 748 8582 800
rect 8754 274 8782 1364
rect 8942 274 8970 1364
rect 9142 872 9148 924
rect 9200 872 9206 924
rect 8736 222 8742 274
rect 8794 222 8800 274
rect 8924 222 8930 274
rect 8982 222 8988 274
rect 9406 150 9434 1364
rect 9538 150 9566 1364
rect 9766 996 9772 1048
rect 9824 996 9830 1048
rect 10002 274 10030 1364
rect 10190 274 10218 1364
rect 10390 1120 10396 1172
rect 10448 1120 10454 1172
rect 9984 222 9990 274
rect 10042 222 10048 274
rect 10172 222 10178 274
rect 10230 222 10236 274
rect 10654 150 10682 1364
rect 10786 150 10814 1364
rect 11014 1244 11020 1296
rect 11072 1244 11078 1296
rect 11250 274 11278 1364
rect 11438 274 11466 1364
rect 11638 376 11644 428
rect 11696 376 11702 428
rect 11232 222 11238 274
rect 11290 222 11296 274
rect 11420 222 11426 274
rect 11478 222 11484 274
rect 11902 150 11930 1364
rect 12034 150 12062 1364
rect 12262 500 12268 552
rect 12320 500 12326 552
rect 12498 274 12526 1364
rect 12686 274 12714 1364
rect 12886 624 12892 676
rect 12944 624 12950 676
rect 12480 222 12486 274
rect 12538 222 12544 274
rect 12668 222 12674 274
rect 12726 222 12732 274
rect 13150 150 13178 1364
rect 13282 150 13310 1364
rect 13510 748 13516 800
rect 13568 748 13574 800
rect 13746 274 13774 1364
rect 13934 274 13962 1364
rect 14134 872 14140 924
rect 14192 872 14198 924
rect 13728 222 13734 274
rect 13786 222 13792 274
rect 13916 222 13922 274
rect 13974 222 13980 274
rect 14398 150 14426 1364
rect 14530 150 14558 1364
rect 14758 996 14764 1048
rect 14816 996 14822 1048
rect 14994 274 15022 1364
rect 15182 274 15210 1364
rect 15382 1120 15388 1172
rect 15440 1120 15446 1172
rect 14976 222 14982 274
rect 15034 222 15040 274
rect 15164 222 15170 274
rect 15222 222 15228 274
rect 15646 150 15674 1364
rect 15778 150 15806 1364
rect 16006 1244 16012 1296
rect 16064 1244 16070 1296
rect 16242 274 16270 1364
rect 16430 274 16458 1364
rect 16630 376 16636 428
rect 16688 376 16694 428
rect 16224 222 16230 274
rect 16282 222 16288 274
rect 16412 222 16418 274
rect 16470 222 16476 274
rect 16894 150 16922 1364
rect 17026 150 17054 1364
rect 17254 500 17260 552
rect 17312 500 17318 552
rect 17490 274 17518 1364
rect 17678 274 17706 1364
rect 17878 624 17884 676
rect 17936 624 17942 676
rect 17472 222 17478 274
rect 17530 222 17536 274
rect 17660 222 17666 274
rect 17718 222 17724 274
rect 18142 150 18170 1364
rect 18274 150 18302 1364
rect 18502 748 18508 800
rect 18560 748 18566 800
rect 18738 274 18766 1364
rect 18926 274 18954 1364
rect 19126 872 19132 924
rect 19184 872 19190 924
rect 18720 222 18726 274
rect 18778 222 18784 274
rect 18908 222 18914 274
rect 18966 222 18972 274
rect 19390 150 19418 1364
rect 19522 150 19550 1364
rect 19750 996 19756 1048
rect 19808 996 19814 1048
rect 19986 274 20014 1364
rect 20174 274 20202 1364
rect 20374 1120 20380 1172
rect 20432 1120 20438 1172
rect 19968 222 19974 274
rect 20026 222 20032 274
rect 20156 222 20162 274
rect 20214 222 20220 274
rect 20638 150 20666 1364
rect 20770 150 20798 1364
rect 20998 1244 21004 1296
rect 21056 1244 21062 1296
rect 21234 274 21262 1364
rect 21422 274 21450 1364
rect 21622 376 21628 428
rect 21680 376 21686 428
rect 21216 222 21222 274
rect 21274 222 21280 274
rect 21404 222 21410 274
rect 21462 222 21468 274
rect 21886 150 21914 1364
rect 22018 150 22046 1364
rect 22246 500 22252 552
rect 22304 500 22310 552
rect 22482 274 22510 1364
rect 22670 274 22698 1364
rect 22870 624 22876 676
rect 22928 624 22934 676
rect 22464 222 22470 274
rect 22522 222 22528 274
rect 22652 222 22658 274
rect 22710 222 22716 274
rect 23134 150 23162 1364
rect 23266 150 23294 1364
rect 23494 748 23500 800
rect 23552 748 23558 800
rect 23730 274 23758 1364
rect 23918 274 23946 1364
rect 24118 872 24124 924
rect 24176 872 24182 924
rect 23712 222 23718 274
rect 23770 222 23776 274
rect 23900 222 23906 274
rect 23958 222 23964 274
rect 24382 150 24410 1364
rect 24514 150 24542 1364
rect 24742 996 24748 1048
rect 24800 996 24806 1048
rect 24978 274 25006 1364
rect 25166 274 25194 1364
rect 25366 1120 25372 1172
rect 25424 1120 25430 1172
rect 24960 222 24966 274
rect 25018 222 25024 274
rect 25148 222 25154 274
rect 25206 222 25212 274
rect 25630 150 25658 1364
rect 25762 150 25790 1364
rect 25990 1244 25996 1296
rect 26048 1244 26054 1296
rect 26226 274 26254 1364
rect 26414 274 26442 1364
rect 26614 376 26620 428
rect 26672 376 26678 428
rect 26208 222 26214 274
rect 26266 222 26272 274
rect 26396 222 26402 274
rect 26454 222 26460 274
rect 26878 150 26906 1364
rect 27010 150 27038 1364
rect 27238 500 27244 552
rect 27296 500 27302 552
rect 27474 274 27502 1364
rect 27662 274 27690 1364
rect 27862 624 27868 676
rect 27920 624 27926 676
rect 27456 222 27462 274
rect 27514 222 27520 274
rect 27644 222 27650 274
rect 27702 222 27708 274
rect 28126 150 28154 1364
rect 28258 150 28286 1364
rect 28486 748 28492 800
rect 28544 748 28550 800
rect 28722 274 28750 1364
rect 28910 274 28938 1364
rect 29110 872 29116 924
rect 29168 872 29174 924
rect 28704 222 28710 274
rect 28762 222 28768 274
rect 28892 222 28898 274
rect 28950 222 28956 274
rect 29374 150 29402 1364
rect 29506 150 29534 1364
rect 29734 996 29740 1048
rect 29792 996 29798 1048
rect 29970 274 29998 1364
rect 30158 274 30186 1364
rect 30358 1120 30364 1172
rect 30416 1120 30422 1172
rect 29952 222 29958 274
rect 30010 222 30016 274
rect 30140 222 30146 274
rect 30198 222 30204 274
rect 30622 150 30650 1364
rect 30754 150 30782 1364
rect 30982 1244 30988 1296
rect 31040 1244 31046 1296
rect 31218 274 31246 1364
rect 31406 274 31434 1364
rect 31606 376 31612 428
rect 31664 376 31670 428
rect 31200 222 31206 274
rect 31258 222 31264 274
rect 31388 222 31394 274
rect 31446 222 31452 274
rect 31870 150 31898 1364
rect 32002 150 32030 1364
rect 32230 500 32236 552
rect 32288 500 32294 552
rect 32466 274 32494 1364
rect 32654 274 32682 1364
rect 32854 624 32860 676
rect 32912 624 32918 676
rect 32448 222 32454 274
rect 32506 222 32512 274
rect 32636 222 32642 274
rect 32694 222 32700 274
rect 33118 150 33146 1364
rect 33250 150 33278 1364
rect 33478 748 33484 800
rect 33536 748 33542 800
rect 33714 274 33742 1364
rect 33902 274 33930 1364
rect 34102 872 34108 924
rect 34160 872 34166 924
rect 33696 222 33702 274
rect 33754 222 33760 274
rect 33884 222 33890 274
rect 33942 222 33948 274
rect 34366 150 34394 1364
rect 34498 150 34526 1364
rect 34726 996 34732 1048
rect 34784 996 34790 1048
rect 34962 274 34990 1364
rect 35150 274 35178 1364
rect 35350 1120 35356 1172
rect 35408 1120 35414 1172
rect 34944 222 34950 274
rect 35002 222 35008 274
rect 35132 222 35138 274
rect 35190 222 35196 274
rect 35614 150 35642 1364
rect 35746 150 35774 1364
rect 35974 1244 35980 1296
rect 36032 1244 36038 1296
rect 36210 274 36238 1364
rect 36398 274 36426 1364
rect 36598 376 36604 428
rect 36656 376 36662 428
rect 36192 222 36198 274
rect 36250 222 36256 274
rect 36380 222 36386 274
rect 36438 222 36444 274
rect 36862 150 36890 1364
rect 36994 150 37022 1364
rect 37222 500 37228 552
rect 37280 500 37286 552
rect 37458 274 37486 1364
rect 37646 274 37674 1364
rect 37846 624 37852 676
rect 37904 624 37910 676
rect 37440 222 37446 274
rect 37498 222 37504 274
rect 37628 222 37634 274
rect 37686 222 37692 274
rect 38110 150 38138 1364
rect 38242 150 38270 1364
rect 38470 748 38476 800
rect 38528 748 38534 800
rect 38706 274 38734 1364
rect 38894 274 38922 1364
rect 39094 872 39100 924
rect 39152 872 39158 924
rect 38688 222 38694 274
rect 38746 222 38752 274
rect 38876 222 38882 274
rect 38934 222 38940 274
rect 39358 150 39386 1364
rect 39490 150 39518 1364
rect 39718 996 39724 1048
rect 39776 996 39782 1048
rect 39954 274 39982 1364
rect 40142 274 40170 1364
rect 40342 1120 40348 1172
rect 40400 1120 40406 1172
rect 39936 222 39942 274
rect 39994 222 40000 274
rect 40124 222 40130 274
rect 40182 222 40188 274
rect 40606 150 40634 1364
rect 40738 150 40766 1364
rect 40966 1244 40972 1296
rect 41024 1244 41030 1296
rect 41202 274 41230 1364
rect 41184 222 41190 274
rect 41242 222 41248 274
rect 1900 98 1906 150
rect 1958 98 1964 150
rect 2032 98 2038 150
rect 2090 98 2096 150
rect 3148 98 3154 150
rect 3206 98 3212 150
rect 3280 98 3286 150
rect 3338 98 3344 150
rect 4396 98 4402 150
rect 4454 98 4460 150
rect 4528 98 4534 150
rect 4586 98 4592 150
rect 5644 98 5650 150
rect 5702 98 5708 150
rect 5776 98 5782 150
rect 5834 98 5840 150
rect 6892 98 6898 150
rect 6950 98 6956 150
rect 7024 98 7030 150
rect 7082 98 7088 150
rect 8140 98 8146 150
rect 8198 98 8204 150
rect 8272 98 8278 150
rect 8330 98 8336 150
rect 9388 98 9394 150
rect 9446 98 9452 150
rect 9520 98 9526 150
rect 9578 98 9584 150
rect 10636 98 10642 150
rect 10694 98 10700 150
rect 10768 98 10774 150
rect 10826 98 10832 150
rect 11884 98 11890 150
rect 11942 98 11948 150
rect 12016 98 12022 150
rect 12074 98 12080 150
rect 13132 98 13138 150
rect 13190 98 13196 150
rect 13264 98 13270 150
rect 13322 98 13328 150
rect 14380 98 14386 150
rect 14438 98 14444 150
rect 14512 98 14518 150
rect 14570 98 14576 150
rect 15628 98 15634 150
rect 15686 98 15692 150
rect 15760 98 15766 150
rect 15818 98 15824 150
rect 16876 98 16882 150
rect 16934 98 16940 150
rect 17008 98 17014 150
rect 17066 98 17072 150
rect 18124 98 18130 150
rect 18182 98 18188 150
rect 18256 98 18262 150
rect 18314 98 18320 150
rect 19372 98 19378 150
rect 19430 98 19436 150
rect 19504 98 19510 150
rect 19562 98 19568 150
rect 20620 98 20626 150
rect 20678 98 20684 150
rect 20752 98 20758 150
rect 20810 98 20816 150
rect 21868 98 21874 150
rect 21926 98 21932 150
rect 22000 98 22006 150
rect 22058 98 22064 150
rect 23116 98 23122 150
rect 23174 98 23180 150
rect 23248 98 23254 150
rect 23306 98 23312 150
rect 24364 98 24370 150
rect 24422 98 24428 150
rect 24496 98 24502 150
rect 24554 98 24560 150
rect 25612 98 25618 150
rect 25670 98 25676 150
rect 25744 98 25750 150
rect 25802 98 25808 150
rect 26860 98 26866 150
rect 26918 98 26924 150
rect 26992 98 26998 150
rect 27050 98 27056 150
rect 28108 98 28114 150
rect 28166 98 28172 150
rect 28240 98 28246 150
rect 28298 98 28304 150
rect 29356 98 29362 150
rect 29414 98 29420 150
rect 29488 98 29494 150
rect 29546 98 29552 150
rect 30604 98 30610 150
rect 30662 98 30668 150
rect 30736 98 30742 150
rect 30794 98 30800 150
rect 31852 98 31858 150
rect 31910 98 31916 150
rect 31984 98 31990 150
rect 32042 98 32048 150
rect 33100 98 33106 150
rect 33158 98 33164 150
rect 33232 98 33238 150
rect 33290 98 33296 150
rect 34348 98 34354 150
rect 34406 98 34412 150
rect 34480 98 34486 150
rect 34538 98 34544 150
rect 35596 98 35602 150
rect 35654 98 35660 150
rect 35728 98 35734 150
rect 35786 98 35792 150
rect 36844 98 36850 150
rect 36902 98 36908 150
rect 36976 98 36982 150
rect 37034 98 37040 150
rect 38092 98 38098 150
rect 38150 98 38156 150
rect 38224 98 38230 150
rect 38282 98 38288 150
rect 39340 98 39346 150
rect 39398 98 39404 150
rect 39472 98 39478 150
rect 39530 98 39536 150
rect 40588 98 40594 150
rect 40646 98 40652 150
rect 40720 98 40726 150
rect 40778 98 40784 150
<< via1 >>
rect 1660 419 1712 428
rect 1660 385 1669 419
rect 1669 385 1703 419
rect 1703 385 1712 419
rect 1660 376 1712 385
rect 1442 222 1494 274
rect 2284 543 2336 552
rect 2284 509 2293 543
rect 2293 509 2327 543
rect 2327 509 2336 543
rect 2284 500 2336 509
rect 2908 667 2960 676
rect 2908 633 2917 667
rect 2917 633 2951 667
rect 2951 633 2960 667
rect 2908 624 2960 633
rect 2502 222 2554 274
rect 2690 222 2742 274
rect 3532 791 3584 800
rect 3532 757 3541 791
rect 3541 757 3575 791
rect 3575 757 3584 791
rect 3532 748 3584 757
rect 4156 915 4208 924
rect 4156 881 4165 915
rect 4165 881 4199 915
rect 4199 881 4208 915
rect 4156 872 4208 881
rect 3750 222 3802 274
rect 3938 222 3990 274
rect 4780 1039 4832 1048
rect 4780 1005 4789 1039
rect 4789 1005 4823 1039
rect 4823 1005 4832 1039
rect 4780 996 4832 1005
rect 5404 1163 5456 1172
rect 5404 1129 5413 1163
rect 5413 1129 5447 1163
rect 5447 1129 5456 1163
rect 5404 1120 5456 1129
rect 4998 222 5050 274
rect 5186 222 5238 274
rect 6028 1287 6080 1296
rect 6028 1253 6037 1287
rect 6037 1253 6071 1287
rect 6071 1253 6080 1287
rect 6028 1244 6080 1253
rect 6652 419 6704 428
rect 6652 385 6661 419
rect 6661 385 6695 419
rect 6695 385 6704 419
rect 6652 376 6704 385
rect 6246 222 6298 274
rect 6434 222 6486 274
rect 7276 543 7328 552
rect 7276 509 7285 543
rect 7285 509 7319 543
rect 7319 509 7328 543
rect 7276 500 7328 509
rect 7900 667 7952 676
rect 7900 633 7909 667
rect 7909 633 7943 667
rect 7943 633 7952 667
rect 7900 624 7952 633
rect 7494 222 7546 274
rect 7682 222 7734 274
rect 8524 791 8576 800
rect 8524 757 8533 791
rect 8533 757 8567 791
rect 8567 757 8576 791
rect 8524 748 8576 757
rect 9148 915 9200 924
rect 9148 881 9157 915
rect 9157 881 9191 915
rect 9191 881 9200 915
rect 9148 872 9200 881
rect 8742 222 8794 274
rect 8930 222 8982 274
rect 9772 1039 9824 1048
rect 9772 1005 9781 1039
rect 9781 1005 9815 1039
rect 9815 1005 9824 1039
rect 9772 996 9824 1005
rect 10396 1163 10448 1172
rect 10396 1129 10405 1163
rect 10405 1129 10439 1163
rect 10439 1129 10448 1163
rect 10396 1120 10448 1129
rect 9990 222 10042 274
rect 10178 222 10230 274
rect 11020 1287 11072 1296
rect 11020 1253 11029 1287
rect 11029 1253 11063 1287
rect 11063 1253 11072 1287
rect 11020 1244 11072 1253
rect 11644 419 11696 428
rect 11644 385 11653 419
rect 11653 385 11687 419
rect 11687 385 11696 419
rect 11644 376 11696 385
rect 11238 222 11290 274
rect 11426 222 11478 274
rect 12268 543 12320 552
rect 12268 509 12277 543
rect 12277 509 12311 543
rect 12311 509 12320 543
rect 12268 500 12320 509
rect 12892 667 12944 676
rect 12892 633 12901 667
rect 12901 633 12935 667
rect 12935 633 12944 667
rect 12892 624 12944 633
rect 12486 222 12538 274
rect 12674 222 12726 274
rect 13516 791 13568 800
rect 13516 757 13525 791
rect 13525 757 13559 791
rect 13559 757 13568 791
rect 13516 748 13568 757
rect 14140 915 14192 924
rect 14140 881 14149 915
rect 14149 881 14183 915
rect 14183 881 14192 915
rect 14140 872 14192 881
rect 13734 222 13786 274
rect 13922 222 13974 274
rect 14764 1039 14816 1048
rect 14764 1005 14773 1039
rect 14773 1005 14807 1039
rect 14807 1005 14816 1039
rect 14764 996 14816 1005
rect 15388 1163 15440 1172
rect 15388 1129 15397 1163
rect 15397 1129 15431 1163
rect 15431 1129 15440 1163
rect 15388 1120 15440 1129
rect 14982 222 15034 274
rect 15170 222 15222 274
rect 16012 1287 16064 1296
rect 16012 1253 16021 1287
rect 16021 1253 16055 1287
rect 16055 1253 16064 1287
rect 16012 1244 16064 1253
rect 16636 419 16688 428
rect 16636 385 16645 419
rect 16645 385 16679 419
rect 16679 385 16688 419
rect 16636 376 16688 385
rect 16230 222 16282 274
rect 16418 222 16470 274
rect 17260 543 17312 552
rect 17260 509 17269 543
rect 17269 509 17303 543
rect 17303 509 17312 543
rect 17260 500 17312 509
rect 17884 667 17936 676
rect 17884 633 17893 667
rect 17893 633 17927 667
rect 17927 633 17936 667
rect 17884 624 17936 633
rect 17478 222 17530 274
rect 17666 222 17718 274
rect 18508 791 18560 800
rect 18508 757 18517 791
rect 18517 757 18551 791
rect 18551 757 18560 791
rect 18508 748 18560 757
rect 19132 915 19184 924
rect 19132 881 19141 915
rect 19141 881 19175 915
rect 19175 881 19184 915
rect 19132 872 19184 881
rect 18726 222 18778 274
rect 18914 222 18966 274
rect 19756 1039 19808 1048
rect 19756 1005 19765 1039
rect 19765 1005 19799 1039
rect 19799 1005 19808 1039
rect 19756 996 19808 1005
rect 20380 1163 20432 1172
rect 20380 1129 20389 1163
rect 20389 1129 20423 1163
rect 20423 1129 20432 1163
rect 20380 1120 20432 1129
rect 19974 222 20026 274
rect 20162 222 20214 274
rect 21004 1287 21056 1296
rect 21004 1253 21013 1287
rect 21013 1253 21047 1287
rect 21047 1253 21056 1287
rect 21004 1244 21056 1253
rect 21628 419 21680 428
rect 21628 385 21637 419
rect 21637 385 21671 419
rect 21671 385 21680 419
rect 21628 376 21680 385
rect 21222 222 21274 274
rect 21410 222 21462 274
rect 22252 543 22304 552
rect 22252 509 22261 543
rect 22261 509 22295 543
rect 22295 509 22304 543
rect 22252 500 22304 509
rect 22876 667 22928 676
rect 22876 633 22885 667
rect 22885 633 22919 667
rect 22919 633 22928 667
rect 22876 624 22928 633
rect 22470 222 22522 274
rect 22658 222 22710 274
rect 23500 791 23552 800
rect 23500 757 23509 791
rect 23509 757 23543 791
rect 23543 757 23552 791
rect 23500 748 23552 757
rect 24124 915 24176 924
rect 24124 881 24133 915
rect 24133 881 24167 915
rect 24167 881 24176 915
rect 24124 872 24176 881
rect 23718 222 23770 274
rect 23906 222 23958 274
rect 24748 1039 24800 1048
rect 24748 1005 24757 1039
rect 24757 1005 24791 1039
rect 24791 1005 24800 1039
rect 24748 996 24800 1005
rect 25372 1163 25424 1172
rect 25372 1129 25381 1163
rect 25381 1129 25415 1163
rect 25415 1129 25424 1163
rect 25372 1120 25424 1129
rect 24966 222 25018 274
rect 25154 222 25206 274
rect 25996 1287 26048 1296
rect 25996 1253 26005 1287
rect 26005 1253 26039 1287
rect 26039 1253 26048 1287
rect 25996 1244 26048 1253
rect 26620 419 26672 428
rect 26620 385 26629 419
rect 26629 385 26663 419
rect 26663 385 26672 419
rect 26620 376 26672 385
rect 26214 222 26266 274
rect 26402 222 26454 274
rect 27244 543 27296 552
rect 27244 509 27253 543
rect 27253 509 27287 543
rect 27287 509 27296 543
rect 27244 500 27296 509
rect 27868 667 27920 676
rect 27868 633 27877 667
rect 27877 633 27911 667
rect 27911 633 27920 667
rect 27868 624 27920 633
rect 27462 222 27514 274
rect 27650 222 27702 274
rect 28492 791 28544 800
rect 28492 757 28501 791
rect 28501 757 28535 791
rect 28535 757 28544 791
rect 28492 748 28544 757
rect 29116 915 29168 924
rect 29116 881 29125 915
rect 29125 881 29159 915
rect 29159 881 29168 915
rect 29116 872 29168 881
rect 28710 222 28762 274
rect 28898 222 28950 274
rect 29740 1039 29792 1048
rect 29740 1005 29749 1039
rect 29749 1005 29783 1039
rect 29783 1005 29792 1039
rect 29740 996 29792 1005
rect 30364 1163 30416 1172
rect 30364 1129 30373 1163
rect 30373 1129 30407 1163
rect 30407 1129 30416 1163
rect 30364 1120 30416 1129
rect 29958 222 30010 274
rect 30146 222 30198 274
rect 30988 1287 31040 1296
rect 30988 1253 30997 1287
rect 30997 1253 31031 1287
rect 31031 1253 31040 1287
rect 30988 1244 31040 1253
rect 31612 419 31664 428
rect 31612 385 31621 419
rect 31621 385 31655 419
rect 31655 385 31664 419
rect 31612 376 31664 385
rect 31206 222 31258 274
rect 31394 222 31446 274
rect 32236 543 32288 552
rect 32236 509 32245 543
rect 32245 509 32279 543
rect 32279 509 32288 543
rect 32236 500 32288 509
rect 32860 667 32912 676
rect 32860 633 32869 667
rect 32869 633 32903 667
rect 32903 633 32912 667
rect 32860 624 32912 633
rect 32454 222 32506 274
rect 32642 222 32694 274
rect 33484 791 33536 800
rect 33484 757 33493 791
rect 33493 757 33527 791
rect 33527 757 33536 791
rect 33484 748 33536 757
rect 34108 915 34160 924
rect 34108 881 34117 915
rect 34117 881 34151 915
rect 34151 881 34160 915
rect 34108 872 34160 881
rect 33702 222 33754 274
rect 33890 222 33942 274
rect 34732 1039 34784 1048
rect 34732 1005 34741 1039
rect 34741 1005 34775 1039
rect 34775 1005 34784 1039
rect 34732 996 34784 1005
rect 35356 1163 35408 1172
rect 35356 1129 35365 1163
rect 35365 1129 35399 1163
rect 35399 1129 35408 1163
rect 35356 1120 35408 1129
rect 34950 222 35002 274
rect 35138 222 35190 274
rect 35980 1287 36032 1296
rect 35980 1253 35989 1287
rect 35989 1253 36023 1287
rect 36023 1253 36032 1287
rect 35980 1244 36032 1253
rect 36604 419 36656 428
rect 36604 385 36613 419
rect 36613 385 36647 419
rect 36647 385 36656 419
rect 36604 376 36656 385
rect 36198 222 36250 274
rect 36386 222 36438 274
rect 37228 543 37280 552
rect 37228 509 37237 543
rect 37237 509 37271 543
rect 37271 509 37280 543
rect 37228 500 37280 509
rect 37852 667 37904 676
rect 37852 633 37861 667
rect 37861 633 37895 667
rect 37895 633 37904 667
rect 37852 624 37904 633
rect 37446 222 37498 274
rect 37634 222 37686 274
rect 38476 791 38528 800
rect 38476 757 38485 791
rect 38485 757 38519 791
rect 38519 757 38528 791
rect 38476 748 38528 757
rect 39100 915 39152 924
rect 39100 881 39109 915
rect 39109 881 39143 915
rect 39143 881 39152 915
rect 39100 872 39152 881
rect 38694 222 38746 274
rect 38882 222 38934 274
rect 39724 1039 39776 1048
rect 39724 1005 39733 1039
rect 39733 1005 39767 1039
rect 39767 1005 39776 1039
rect 39724 996 39776 1005
rect 40348 1163 40400 1172
rect 40348 1129 40357 1163
rect 40357 1129 40391 1163
rect 40391 1129 40400 1163
rect 40348 1120 40400 1129
rect 39942 222 39994 274
rect 40130 222 40182 274
rect 40972 1287 41024 1296
rect 40972 1253 40981 1287
rect 40981 1253 41015 1287
rect 41015 1253 41024 1287
rect 40972 1244 41024 1253
rect 41190 222 41242 274
rect 1906 98 1958 150
rect 2038 98 2090 150
rect 3154 98 3206 150
rect 3286 98 3338 150
rect 4402 98 4454 150
rect 4534 98 4586 150
rect 5650 98 5702 150
rect 5782 98 5834 150
rect 6898 98 6950 150
rect 7030 98 7082 150
rect 8146 98 8198 150
rect 8278 98 8330 150
rect 9394 98 9446 150
rect 9526 98 9578 150
rect 10642 98 10694 150
rect 10774 98 10826 150
rect 11890 98 11942 150
rect 12022 98 12074 150
rect 13138 98 13190 150
rect 13270 98 13322 150
rect 14386 98 14438 150
rect 14518 98 14570 150
rect 15634 98 15686 150
rect 15766 98 15818 150
rect 16882 98 16934 150
rect 17014 98 17066 150
rect 18130 98 18182 150
rect 18262 98 18314 150
rect 19378 98 19430 150
rect 19510 98 19562 150
rect 20626 98 20678 150
rect 20758 98 20810 150
rect 21874 98 21926 150
rect 22006 98 22058 150
rect 23122 98 23174 150
rect 23254 98 23306 150
rect 24370 98 24422 150
rect 24502 98 24554 150
rect 25618 98 25670 150
rect 25750 98 25802 150
rect 26866 98 26918 150
rect 26998 98 27050 150
rect 28114 98 28166 150
rect 28246 98 28298 150
rect 29362 98 29414 150
rect 29494 98 29546 150
rect 30610 98 30662 150
rect 30742 98 30794 150
rect 31858 98 31910 150
rect 31990 98 32042 150
rect 33106 98 33158 150
rect 33238 98 33290 150
rect 34354 98 34406 150
rect 34486 98 34538 150
rect 35602 98 35654 150
rect 35734 98 35786 150
rect 36850 98 36902 150
rect 36982 98 37034 150
rect 38098 98 38150 150
rect 38230 98 38282 150
rect 39346 98 39398 150
rect 39478 98 39530 150
rect 40594 98 40646 150
rect 40726 98 40778 150
<< metal2 >>
rect 6026 1298 6082 1307
rect 6026 1233 6082 1242
rect 11018 1298 11074 1307
rect 11018 1233 11074 1242
rect 16010 1298 16066 1307
rect 16010 1233 16066 1242
rect 21002 1298 21058 1307
rect 21002 1233 21058 1242
rect 25994 1298 26050 1307
rect 25994 1233 26050 1242
rect 30986 1298 31042 1307
rect 30986 1233 31042 1242
rect 35978 1298 36034 1307
rect 35978 1233 36034 1242
rect 40970 1298 41026 1307
rect 40970 1233 41026 1242
rect 5402 1174 5458 1183
rect 5402 1109 5458 1118
rect 10394 1174 10450 1183
rect 10394 1109 10450 1118
rect 15386 1174 15442 1183
rect 15386 1109 15442 1118
rect 20378 1174 20434 1183
rect 20378 1109 20434 1118
rect 25370 1174 25426 1183
rect 25370 1109 25426 1118
rect 30362 1174 30418 1183
rect 30362 1109 30418 1118
rect 35354 1174 35410 1183
rect 35354 1109 35410 1118
rect 40346 1174 40402 1183
rect 40346 1109 40402 1118
rect 4778 1050 4834 1059
rect 4778 985 4834 994
rect 9770 1050 9826 1059
rect 9770 985 9826 994
rect 14762 1050 14818 1059
rect 14762 985 14818 994
rect 19754 1050 19810 1059
rect 19754 985 19810 994
rect 24746 1050 24802 1059
rect 24746 985 24802 994
rect 29738 1050 29794 1059
rect 29738 985 29794 994
rect 34730 1050 34786 1059
rect 34730 985 34786 994
rect 39722 1050 39778 1059
rect 39722 985 39778 994
rect 4154 926 4210 935
rect 4154 861 4210 870
rect 9146 926 9202 935
rect 9146 861 9202 870
rect 14138 926 14194 935
rect 14138 861 14194 870
rect 19130 926 19186 935
rect 19130 861 19186 870
rect 24122 926 24178 935
rect 24122 861 24178 870
rect 29114 926 29170 935
rect 29114 861 29170 870
rect 34106 926 34162 935
rect 34106 861 34162 870
rect 39098 926 39154 935
rect 39098 861 39154 870
rect 3530 802 3586 811
rect 3530 737 3586 746
rect 8522 802 8578 811
rect 8522 737 8578 746
rect 13514 802 13570 811
rect 13514 737 13570 746
rect 18506 802 18562 811
rect 18506 737 18562 746
rect 23498 802 23554 811
rect 23498 737 23554 746
rect 28490 802 28546 811
rect 28490 737 28546 746
rect 33482 802 33538 811
rect 33482 737 33538 746
rect 38474 802 38530 811
rect 38474 737 38530 746
rect 2906 678 2962 687
rect 2906 613 2962 622
rect 7898 678 7954 687
rect 7898 613 7954 622
rect 12890 678 12946 687
rect 12890 613 12946 622
rect 17882 678 17938 687
rect 17882 613 17938 622
rect 22874 678 22930 687
rect 22874 613 22930 622
rect 27866 678 27922 687
rect 27866 613 27922 622
rect 32858 678 32914 687
rect 32858 613 32914 622
rect 37850 678 37906 687
rect 37850 613 37906 622
rect 2282 554 2338 563
rect 2282 489 2338 498
rect 7274 554 7330 563
rect 7274 489 7330 498
rect 12266 554 12322 563
rect 12266 489 12322 498
rect 17258 554 17314 563
rect 17258 489 17314 498
rect 22250 554 22306 563
rect 22250 489 22306 498
rect 27242 554 27298 563
rect 27242 489 27298 498
rect 32234 554 32290 563
rect 32234 489 32290 498
rect 37226 554 37282 563
rect 37226 489 37282 498
rect 1658 430 1714 439
rect 1658 365 1714 374
rect 6650 430 6706 439
rect 6650 365 6706 374
rect 11642 430 11698 439
rect 11642 365 11698 374
rect 16634 430 16690 439
rect 16634 365 16690 374
rect 21626 430 21682 439
rect 21626 365 21682 374
rect 26618 430 26674 439
rect 26618 365 26674 374
rect 31610 430 31666 439
rect 31610 365 31666 374
rect 36602 430 36658 439
rect 36602 365 36658 374
rect 1440 276 1496 285
rect 1440 211 1496 220
rect 2500 276 2556 285
rect 2500 211 2556 220
rect 2688 276 2744 285
rect 2688 211 2744 220
rect 3748 276 3804 285
rect 3748 211 3804 220
rect 3936 276 3992 285
rect 3936 211 3992 220
rect 4996 276 5052 285
rect 4996 211 5052 220
rect 5184 276 5240 285
rect 5184 211 5240 220
rect 6244 276 6300 285
rect 6244 211 6300 220
rect 6432 276 6488 285
rect 6432 211 6488 220
rect 7492 276 7548 285
rect 7492 211 7548 220
rect 7680 276 7736 285
rect 7680 211 7736 220
rect 8740 276 8796 285
rect 8740 211 8796 220
rect 8928 276 8984 285
rect 8928 211 8984 220
rect 9988 276 10044 285
rect 9988 211 10044 220
rect 10176 276 10232 285
rect 10176 211 10232 220
rect 11236 276 11292 285
rect 11236 211 11292 220
rect 11424 276 11480 285
rect 11424 211 11480 220
rect 12484 276 12540 285
rect 12484 211 12540 220
rect 12672 276 12728 285
rect 12672 211 12728 220
rect 13732 276 13788 285
rect 13732 211 13788 220
rect 13920 276 13976 285
rect 13920 211 13976 220
rect 14980 276 15036 285
rect 14980 211 15036 220
rect 15168 276 15224 285
rect 15168 211 15224 220
rect 16228 276 16284 285
rect 16228 211 16284 220
rect 16416 276 16472 285
rect 16416 211 16472 220
rect 17476 276 17532 285
rect 17476 211 17532 220
rect 17664 276 17720 285
rect 17664 211 17720 220
rect 18724 276 18780 285
rect 18724 211 18780 220
rect 18912 276 18968 285
rect 18912 211 18968 220
rect 19972 276 20028 285
rect 19972 211 20028 220
rect 20160 276 20216 285
rect 20160 211 20216 220
rect 21220 276 21276 285
rect 21220 211 21276 220
rect 21408 276 21464 285
rect 21408 211 21464 220
rect 22468 276 22524 285
rect 22468 211 22524 220
rect 22656 276 22712 285
rect 22656 211 22712 220
rect 23716 276 23772 285
rect 23716 211 23772 220
rect 23904 276 23960 285
rect 23904 211 23960 220
rect 24964 276 25020 285
rect 24964 211 25020 220
rect 25152 276 25208 285
rect 25152 211 25208 220
rect 26212 276 26268 285
rect 26212 211 26268 220
rect 26400 276 26456 285
rect 26400 211 26456 220
rect 27460 276 27516 285
rect 27460 211 27516 220
rect 27648 276 27704 285
rect 27648 211 27704 220
rect 28708 276 28764 285
rect 28708 211 28764 220
rect 28896 276 28952 285
rect 28896 211 28952 220
rect 29956 276 30012 285
rect 29956 211 30012 220
rect 30144 276 30200 285
rect 30144 211 30200 220
rect 31204 276 31260 285
rect 31204 211 31260 220
rect 31392 276 31448 285
rect 31392 211 31448 220
rect 32452 276 32508 285
rect 32452 211 32508 220
rect 32640 276 32696 285
rect 32640 211 32696 220
rect 33700 276 33756 285
rect 33700 211 33756 220
rect 33888 276 33944 285
rect 33888 211 33944 220
rect 34948 276 35004 285
rect 34948 211 35004 220
rect 35136 276 35192 285
rect 35136 211 35192 220
rect 36196 276 36252 285
rect 36196 211 36252 220
rect 36384 276 36440 285
rect 36384 211 36440 220
rect 37444 276 37500 285
rect 37444 211 37500 220
rect 37632 276 37688 285
rect 37632 211 37688 220
rect 38692 276 38748 285
rect 38692 211 38748 220
rect 38880 276 38936 285
rect 38880 211 38936 220
rect 39940 276 39996 285
rect 39940 211 39996 220
rect 40128 276 40184 285
rect 40128 211 40184 220
rect 41188 276 41244 285
rect 41188 211 41244 220
rect 1904 152 1960 161
rect 1904 87 1960 96
rect 2036 152 2092 161
rect 2036 87 2092 96
rect 3152 152 3208 161
rect 3152 87 3208 96
rect 3284 152 3340 161
rect 3284 87 3340 96
rect 4400 152 4456 161
rect 4400 87 4456 96
rect 4532 152 4588 161
rect 4532 87 4588 96
rect 5648 152 5704 161
rect 5648 87 5704 96
rect 5780 152 5836 161
rect 5780 87 5836 96
rect 6896 152 6952 161
rect 6896 87 6952 96
rect 7028 152 7084 161
rect 7028 87 7084 96
rect 8144 152 8200 161
rect 8144 87 8200 96
rect 8276 152 8332 161
rect 8276 87 8332 96
rect 9392 152 9448 161
rect 9392 87 9448 96
rect 9524 152 9580 161
rect 9524 87 9580 96
rect 10640 152 10696 161
rect 10640 87 10696 96
rect 10772 152 10828 161
rect 10772 87 10828 96
rect 11888 152 11944 161
rect 11888 87 11944 96
rect 12020 152 12076 161
rect 12020 87 12076 96
rect 13136 152 13192 161
rect 13136 87 13192 96
rect 13268 152 13324 161
rect 13268 87 13324 96
rect 14384 152 14440 161
rect 14384 87 14440 96
rect 14516 152 14572 161
rect 14516 87 14572 96
rect 15632 152 15688 161
rect 15632 87 15688 96
rect 15764 152 15820 161
rect 15764 87 15820 96
rect 16880 152 16936 161
rect 16880 87 16936 96
rect 17012 152 17068 161
rect 17012 87 17068 96
rect 18128 152 18184 161
rect 18128 87 18184 96
rect 18260 152 18316 161
rect 18260 87 18316 96
rect 19376 152 19432 161
rect 19376 87 19432 96
rect 19508 152 19564 161
rect 19508 87 19564 96
rect 20624 152 20680 161
rect 20624 87 20680 96
rect 20756 152 20812 161
rect 20756 87 20812 96
rect 21872 152 21928 161
rect 21872 87 21928 96
rect 22004 152 22060 161
rect 22004 87 22060 96
rect 23120 152 23176 161
rect 23120 87 23176 96
rect 23252 152 23308 161
rect 23252 87 23308 96
rect 24368 152 24424 161
rect 24368 87 24424 96
rect 24500 152 24556 161
rect 24500 87 24556 96
rect 25616 152 25672 161
rect 25616 87 25672 96
rect 25748 152 25804 161
rect 25748 87 25804 96
rect 26864 152 26920 161
rect 26864 87 26920 96
rect 26996 152 27052 161
rect 26996 87 27052 96
rect 28112 152 28168 161
rect 28112 87 28168 96
rect 28244 152 28300 161
rect 28244 87 28300 96
rect 29360 152 29416 161
rect 29360 87 29416 96
rect 29492 152 29548 161
rect 29492 87 29548 96
rect 30608 152 30664 161
rect 30608 87 30664 96
rect 30740 152 30796 161
rect 30740 87 30796 96
rect 31856 152 31912 161
rect 31856 87 31912 96
rect 31988 152 32044 161
rect 31988 87 32044 96
rect 33104 152 33160 161
rect 33104 87 33160 96
rect 33236 152 33292 161
rect 33236 87 33292 96
rect 34352 152 34408 161
rect 34352 87 34408 96
rect 34484 152 34540 161
rect 34484 87 34540 96
rect 35600 152 35656 161
rect 35600 87 35656 96
rect 35732 152 35788 161
rect 35732 87 35788 96
rect 36848 152 36904 161
rect 36848 87 36904 96
rect 36980 152 37036 161
rect 36980 87 37036 96
rect 38096 152 38152 161
rect 38096 87 38152 96
rect 38228 152 38284 161
rect 38228 87 38284 96
rect 39344 152 39400 161
rect 39344 87 39400 96
rect 39476 152 39532 161
rect 39476 87 39532 96
rect 40592 152 40648 161
rect 40592 87 40648 96
rect 40724 152 40780 161
rect 40724 87 40780 96
<< via2 >>
rect 6026 1296 6082 1298
rect 6026 1244 6028 1296
rect 6028 1244 6080 1296
rect 6080 1244 6082 1296
rect 6026 1242 6082 1244
rect 11018 1296 11074 1298
rect 11018 1244 11020 1296
rect 11020 1244 11072 1296
rect 11072 1244 11074 1296
rect 11018 1242 11074 1244
rect 16010 1296 16066 1298
rect 16010 1244 16012 1296
rect 16012 1244 16064 1296
rect 16064 1244 16066 1296
rect 16010 1242 16066 1244
rect 21002 1296 21058 1298
rect 21002 1244 21004 1296
rect 21004 1244 21056 1296
rect 21056 1244 21058 1296
rect 21002 1242 21058 1244
rect 25994 1296 26050 1298
rect 25994 1244 25996 1296
rect 25996 1244 26048 1296
rect 26048 1244 26050 1296
rect 25994 1242 26050 1244
rect 30986 1296 31042 1298
rect 30986 1244 30988 1296
rect 30988 1244 31040 1296
rect 31040 1244 31042 1296
rect 30986 1242 31042 1244
rect 35978 1296 36034 1298
rect 35978 1244 35980 1296
rect 35980 1244 36032 1296
rect 36032 1244 36034 1296
rect 35978 1242 36034 1244
rect 40970 1296 41026 1298
rect 40970 1244 40972 1296
rect 40972 1244 41024 1296
rect 41024 1244 41026 1296
rect 40970 1242 41026 1244
rect 5402 1172 5458 1174
rect 5402 1120 5404 1172
rect 5404 1120 5456 1172
rect 5456 1120 5458 1172
rect 5402 1118 5458 1120
rect 10394 1172 10450 1174
rect 10394 1120 10396 1172
rect 10396 1120 10448 1172
rect 10448 1120 10450 1172
rect 10394 1118 10450 1120
rect 15386 1172 15442 1174
rect 15386 1120 15388 1172
rect 15388 1120 15440 1172
rect 15440 1120 15442 1172
rect 15386 1118 15442 1120
rect 20378 1172 20434 1174
rect 20378 1120 20380 1172
rect 20380 1120 20432 1172
rect 20432 1120 20434 1172
rect 20378 1118 20434 1120
rect 25370 1172 25426 1174
rect 25370 1120 25372 1172
rect 25372 1120 25424 1172
rect 25424 1120 25426 1172
rect 25370 1118 25426 1120
rect 30362 1172 30418 1174
rect 30362 1120 30364 1172
rect 30364 1120 30416 1172
rect 30416 1120 30418 1172
rect 30362 1118 30418 1120
rect 35354 1172 35410 1174
rect 35354 1120 35356 1172
rect 35356 1120 35408 1172
rect 35408 1120 35410 1172
rect 35354 1118 35410 1120
rect 40346 1172 40402 1174
rect 40346 1120 40348 1172
rect 40348 1120 40400 1172
rect 40400 1120 40402 1172
rect 40346 1118 40402 1120
rect 4778 1048 4834 1050
rect 4778 996 4780 1048
rect 4780 996 4832 1048
rect 4832 996 4834 1048
rect 4778 994 4834 996
rect 9770 1048 9826 1050
rect 9770 996 9772 1048
rect 9772 996 9824 1048
rect 9824 996 9826 1048
rect 9770 994 9826 996
rect 14762 1048 14818 1050
rect 14762 996 14764 1048
rect 14764 996 14816 1048
rect 14816 996 14818 1048
rect 14762 994 14818 996
rect 19754 1048 19810 1050
rect 19754 996 19756 1048
rect 19756 996 19808 1048
rect 19808 996 19810 1048
rect 19754 994 19810 996
rect 24746 1048 24802 1050
rect 24746 996 24748 1048
rect 24748 996 24800 1048
rect 24800 996 24802 1048
rect 24746 994 24802 996
rect 29738 1048 29794 1050
rect 29738 996 29740 1048
rect 29740 996 29792 1048
rect 29792 996 29794 1048
rect 29738 994 29794 996
rect 34730 1048 34786 1050
rect 34730 996 34732 1048
rect 34732 996 34784 1048
rect 34784 996 34786 1048
rect 34730 994 34786 996
rect 39722 1048 39778 1050
rect 39722 996 39724 1048
rect 39724 996 39776 1048
rect 39776 996 39778 1048
rect 39722 994 39778 996
rect 4154 924 4210 926
rect 4154 872 4156 924
rect 4156 872 4208 924
rect 4208 872 4210 924
rect 4154 870 4210 872
rect 9146 924 9202 926
rect 9146 872 9148 924
rect 9148 872 9200 924
rect 9200 872 9202 924
rect 9146 870 9202 872
rect 14138 924 14194 926
rect 14138 872 14140 924
rect 14140 872 14192 924
rect 14192 872 14194 924
rect 14138 870 14194 872
rect 19130 924 19186 926
rect 19130 872 19132 924
rect 19132 872 19184 924
rect 19184 872 19186 924
rect 19130 870 19186 872
rect 24122 924 24178 926
rect 24122 872 24124 924
rect 24124 872 24176 924
rect 24176 872 24178 924
rect 24122 870 24178 872
rect 29114 924 29170 926
rect 29114 872 29116 924
rect 29116 872 29168 924
rect 29168 872 29170 924
rect 29114 870 29170 872
rect 34106 924 34162 926
rect 34106 872 34108 924
rect 34108 872 34160 924
rect 34160 872 34162 924
rect 34106 870 34162 872
rect 39098 924 39154 926
rect 39098 872 39100 924
rect 39100 872 39152 924
rect 39152 872 39154 924
rect 39098 870 39154 872
rect 3530 800 3586 802
rect 3530 748 3532 800
rect 3532 748 3584 800
rect 3584 748 3586 800
rect 3530 746 3586 748
rect 8522 800 8578 802
rect 8522 748 8524 800
rect 8524 748 8576 800
rect 8576 748 8578 800
rect 8522 746 8578 748
rect 13514 800 13570 802
rect 13514 748 13516 800
rect 13516 748 13568 800
rect 13568 748 13570 800
rect 13514 746 13570 748
rect 18506 800 18562 802
rect 18506 748 18508 800
rect 18508 748 18560 800
rect 18560 748 18562 800
rect 18506 746 18562 748
rect 23498 800 23554 802
rect 23498 748 23500 800
rect 23500 748 23552 800
rect 23552 748 23554 800
rect 23498 746 23554 748
rect 28490 800 28546 802
rect 28490 748 28492 800
rect 28492 748 28544 800
rect 28544 748 28546 800
rect 28490 746 28546 748
rect 33482 800 33538 802
rect 33482 748 33484 800
rect 33484 748 33536 800
rect 33536 748 33538 800
rect 33482 746 33538 748
rect 38474 800 38530 802
rect 38474 748 38476 800
rect 38476 748 38528 800
rect 38528 748 38530 800
rect 38474 746 38530 748
rect 2906 676 2962 678
rect 2906 624 2908 676
rect 2908 624 2960 676
rect 2960 624 2962 676
rect 2906 622 2962 624
rect 7898 676 7954 678
rect 7898 624 7900 676
rect 7900 624 7952 676
rect 7952 624 7954 676
rect 7898 622 7954 624
rect 12890 676 12946 678
rect 12890 624 12892 676
rect 12892 624 12944 676
rect 12944 624 12946 676
rect 12890 622 12946 624
rect 17882 676 17938 678
rect 17882 624 17884 676
rect 17884 624 17936 676
rect 17936 624 17938 676
rect 17882 622 17938 624
rect 22874 676 22930 678
rect 22874 624 22876 676
rect 22876 624 22928 676
rect 22928 624 22930 676
rect 22874 622 22930 624
rect 27866 676 27922 678
rect 27866 624 27868 676
rect 27868 624 27920 676
rect 27920 624 27922 676
rect 27866 622 27922 624
rect 32858 676 32914 678
rect 32858 624 32860 676
rect 32860 624 32912 676
rect 32912 624 32914 676
rect 32858 622 32914 624
rect 37850 676 37906 678
rect 37850 624 37852 676
rect 37852 624 37904 676
rect 37904 624 37906 676
rect 37850 622 37906 624
rect 2282 552 2338 554
rect 2282 500 2284 552
rect 2284 500 2336 552
rect 2336 500 2338 552
rect 2282 498 2338 500
rect 7274 552 7330 554
rect 7274 500 7276 552
rect 7276 500 7328 552
rect 7328 500 7330 552
rect 7274 498 7330 500
rect 12266 552 12322 554
rect 12266 500 12268 552
rect 12268 500 12320 552
rect 12320 500 12322 552
rect 12266 498 12322 500
rect 17258 552 17314 554
rect 17258 500 17260 552
rect 17260 500 17312 552
rect 17312 500 17314 552
rect 17258 498 17314 500
rect 22250 552 22306 554
rect 22250 500 22252 552
rect 22252 500 22304 552
rect 22304 500 22306 552
rect 22250 498 22306 500
rect 27242 552 27298 554
rect 27242 500 27244 552
rect 27244 500 27296 552
rect 27296 500 27298 552
rect 27242 498 27298 500
rect 32234 552 32290 554
rect 32234 500 32236 552
rect 32236 500 32288 552
rect 32288 500 32290 552
rect 32234 498 32290 500
rect 37226 552 37282 554
rect 37226 500 37228 552
rect 37228 500 37280 552
rect 37280 500 37282 552
rect 37226 498 37282 500
rect 1658 428 1714 430
rect 1658 376 1660 428
rect 1660 376 1712 428
rect 1712 376 1714 428
rect 1658 374 1714 376
rect 6650 428 6706 430
rect 6650 376 6652 428
rect 6652 376 6704 428
rect 6704 376 6706 428
rect 6650 374 6706 376
rect 11642 428 11698 430
rect 11642 376 11644 428
rect 11644 376 11696 428
rect 11696 376 11698 428
rect 11642 374 11698 376
rect 16634 428 16690 430
rect 16634 376 16636 428
rect 16636 376 16688 428
rect 16688 376 16690 428
rect 16634 374 16690 376
rect 21626 428 21682 430
rect 21626 376 21628 428
rect 21628 376 21680 428
rect 21680 376 21682 428
rect 21626 374 21682 376
rect 26618 428 26674 430
rect 26618 376 26620 428
rect 26620 376 26672 428
rect 26672 376 26674 428
rect 26618 374 26674 376
rect 31610 428 31666 430
rect 31610 376 31612 428
rect 31612 376 31664 428
rect 31664 376 31666 428
rect 31610 374 31666 376
rect 36602 428 36658 430
rect 36602 376 36604 428
rect 36604 376 36656 428
rect 36656 376 36658 428
rect 36602 374 36658 376
rect 1440 274 1496 276
rect 1440 222 1442 274
rect 1442 222 1494 274
rect 1494 222 1496 274
rect 1440 220 1496 222
rect 2500 274 2556 276
rect 2500 222 2502 274
rect 2502 222 2554 274
rect 2554 222 2556 274
rect 2500 220 2556 222
rect 2688 274 2744 276
rect 2688 222 2690 274
rect 2690 222 2742 274
rect 2742 222 2744 274
rect 2688 220 2744 222
rect 3748 274 3804 276
rect 3748 222 3750 274
rect 3750 222 3802 274
rect 3802 222 3804 274
rect 3748 220 3804 222
rect 3936 274 3992 276
rect 3936 222 3938 274
rect 3938 222 3990 274
rect 3990 222 3992 274
rect 3936 220 3992 222
rect 4996 274 5052 276
rect 4996 222 4998 274
rect 4998 222 5050 274
rect 5050 222 5052 274
rect 4996 220 5052 222
rect 5184 274 5240 276
rect 5184 222 5186 274
rect 5186 222 5238 274
rect 5238 222 5240 274
rect 5184 220 5240 222
rect 6244 274 6300 276
rect 6244 222 6246 274
rect 6246 222 6298 274
rect 6298 222 6300 274
rect 6244 220 6300 222
rect 6432 274 6488 276
rect 6432 222 6434 274
rect 6434 222 6486 274
rect 6486 222 6488 274
rect 6432 220 6488 222
rect 7492 274 7548 276
rect 7492 222 7494 274
rect 7494 222 7546 274
rect 7546 222 7548 274
rect 7492 220 7548 222
rect 7680 274 7736 276
rect 7680 222 7682 274
rect 7682 222 7734 274
rect 7734 222 7736 274
rect 7680 220 7736 222
rect 8740 274 8796 276
rect 8740 222 8742 274
rect 8742 222 8794 274
rect 8794 222 8796 274
rect 8740 220 8796 222
rect 8928 274 8984 276
rect 8928 222 8930 274
rect 8930 222 8982 274
rect 8982 222 8984 274
rect 8928 220 8984 222
rect 9988 274 10044 276
rect 9988 222 9990 274
rect 9990 222 10042 274
rect 10042 222 10044 274
rect 9988 220 10044 222
rect 10176 274 10232 276
rect 10176 222 10178 274
rect 10178 222 10230 274
rect 10230 222 10232 274
rect 10176 220 10232 222
rect 11236 274 11292 276
rect 11236 222 11238 274
rect 11238 222 11290 274
rect 11290 222 11292 274
rect 11236 220 11292 222
rect 11424 274 11480 276
rect 11424 222 11426 274
rect 11426 222 11478 274
rect 11478 222 11480 274
rect 11424 220 11480 222
rect 12484 274 12540 276
rect 12484 222 12486 274
rect 12486 222 12538 274
rect 12538 222 12540 274
rect 12484 220 12540 222
rect 12672 274 12728 276
rect 12672 222 12674 274
rect 12674 222 12726 274
rect 12726 222 12728 274
rect 12672 220 12728 222
rect 13732 274 13788 276
rect 13732 222 13734 274
rect 13734 222 13786 274
rect 13786 222 13788 274
rect 13732 220 13788 222
rect 13920 274 13976 276
rect 13920 222 13922 274
rect 13922 222 13974 274
rect 13974 222 13976 274
rect 13920 220 13976 222
rect 14980 274 15036 276
rect 14980 222 14982 274
rect 14982 222 15034 274
rect 15034 222 15036 274
rect 14980 220 15036 222
rect 15168 274 15224 276
rect 15168 222 15170 274
rect 15170 222 15222 274
rect 15222 222 15224 274
rect 15168 220 15224 222
rect 16228 274 16284 276
rect 16228 222 16230 274
rect 16230 222 16282 274
rect 16282 222 16284 274
rect 16228 220 16284 222
rect 16416 274 16472 276
rect 16416 222 16418 274
rect 16418 222 16470 274
rect 16470 222 16472 274
rect 16416 220 16472 222
rect 17476 274 17532 276
rect 17476 222 17478 274
rect 17478 222 17530 274
rect 17530 222 17532 274
rect 17476 220 17532 222
rect 17664 274 17720 276
rect 17664 222 17666 274
rect 17666 222 17718 274
rect 17718 222 17720 274
rect 17664 220 17720 222
rect 18724 274 18780 276
rect 18724 222 18726 274
rect 18726 222 18778 274
rect 18778 222 18780 274
rect 18724 220 18780 222
rect 18912 274 18968 276
rect 18912 222 18914 274
rect 18914 222 18966 274
rect 18966 222 18968 274
rect 18912 220 18968 222
rect 19972 274 20028 276
rect 19972 222 19974 274
rect 19974 222 20026 274
rect 20026 222 20028 274
rect 19972 220 20028 222
rect 20160 274 20216 276
rect 20160 222 20162 274
rect 20162 222 20214 274
rect 20214 222 20216 274
rect 20160 220 20216 222
rect 21220 274 21276 276
rect 21220 222 21222 274
rect 21222 222 21274 274
rect 21274 222 21276 274
rect 21220 220 21276 222
rect 21408 274 21464 276
rect 21408 222 21410 274
rect 21410 222 21462 274
rect 21462 222 21464 274
rect 21408 220 21464 222
rect 22468 274 22524 276
rect 22468 222 22470 274
rect 22470 222 22522 274
rect 22522 222 22524 274
rect 22468 220 22524 222
rect 22656 274 22712 276
rect 22656 222 22658 274
rect 22658 222 22710 274
rect 22710 222 22712 274
rect 22656 220 22712 222
rect 23716 274 23772 276
rect 23716 222 23718 274
rect 23718 222 23770 274
rect 23770 222 23772 274
rect 23716 220 23772 222
rect 23904 274 23960 276
rect 23904 222 23906 274
rect 23906 222 23958 274
rect 23958 222 23960 274
rect 23904 220 23960 222
rect 24964 274 25020 276
rect 24964 222 24966 274
rect 24966 222 25018 274
rect 25018 222 25020 274
rect 24964 220 25020 222
rect 25152 274 25208 276
rect 25152 222 25154 274
rect 25154 222 25206 274
rect 25206 222 25208 274
rect 25152 220 25208 222
rect 26212 274 26268 276
rect 26212 222 26214 274
rect 26214 222 26266 274
rect 26266 222 26268 274
rect 26212 220 26268 222
rect 26400 274 26456 276
rect 26400 222 26402 274
rect 26402 222 26454 274
rect 26454 222 26456 274
rect 26400 220 26456 222
rect 27460 274 27516 276
rect 27460 222 27462 274
rect 27462 222 27514 274
rect 27514 222 27516 274
rect 27460 220 27516 222
rect 27648 274 27704 276
rect 27648 222 27650 274
rect 27650 222 27702 274
rect 27702 222 27704 274
rect 27648 220 27704 222
rect 28708 274 28764 276
rect 28708 222 28710 274
rect 28710 222 28762 274
rect 28762 222 28764 274
rect 28708 220 28764 222
rect 28896 274 28952 276
rect 28896 222 28898 274
rect 28898 222 28950 274
rect 28950 222 28952 274
rect 28896 220 28952 222
rect 29956 274 30012 276
rect 29956 222 29958 274
rect 29958 222 30010 274
rect 30010 222 30012 274
rect 29956 220 30012 222
rect 30144 274 30200 276
rect 30144 222 30146 274
rect 30146 222 30198 274
rect 30198 222 30200 274
rect 30144 220 30200 222
rect 31204 274 31260 276
rect 31204 222 31206 274
rect 31206 222 31258 274
rect 31258 222 31260 274
rect 31204 220 31260 222
rect 31392 274 31448 276
rect 31392 222 31394 274
rect 31394 222 31446 274
rect 31446 222 31448 274
rect 31392 220 31448 222
rect 32452 274 32508 276
rect 32452 222 32454 274
rect 32454 222 32506 274
rect 32506 222 32508 274
rect 32452 220 32508 222
rect 32640 274 32696 276
rect 32640 222 32642 274
rect 32642 222 32694 274
rect 32694 222 32696 274
rect 32640 220 32696 222
rect 33700 274 33756 276
rect 33700 222 33702 274
rect 33702 222 33754 274
rect 33754 222 33756 274
rect 33700 220 33756 222
rect 33888 274 33944 276
rect 33888 222 33890 274
rect 33890 222 33942 274
rect 33942 222 33944 274
rect 33888 220 33944 222
rect 34948 274 35004 276
rect 34948 222 34950 274
rect 34950 222 35002 274
rect 35002 222 35004 274
rect 34948 220 35004 222
rect 35136 274 35192 276
rect 35136 222 35138 274
rect 35138 222 35190 274
rect 35190 222 35192 274
rect 35136 220 35192 222
rect 36196 274 36252 276
rect 36196 222 36198 274
rect 36198 222 36250 274
rect 36250 222 36252 274
rect 36196 220 36252 222
rect 36384 274 36440 276
rect 36384 222 36386 274
rect 36386 222 36438 274
rect 36438 222 36440 274
rect 36384 220 36440 222
rect 37444 274 37500 276
rect 37444 222 37446 274
rect 37446 222 37498 274
rect 37498 222 37500 274
rect 37444 220 37500 222
rect 37632 274 37688 276
rect 37632 222 37634 274
rect 37634 222 37686 274
rect 37686 222 37688 274
rect 37632 220 37688 222
rect 38692 274 38748 276
rect 38692 222 38694 274
rect 38694 222 38746 274
rect 38746 222 38748 274
rect 38692 220 38748 222
rect 38880 274 38936 276
rect 38880 222 38882 274
rect 38882 222 38934 274
rect 38934 222 38936 274
rect 38880 220 38936 222
rect 39940 274 39996 276
rect 39940 222 39942 274
rect 39942 222 39994 274
rect 39994 222 39996 274
rect 39940 220 39996 222
rect 40128 274 40184 276
rect 40128 222 40130 274
rect 40130 222 40182 274
rect 40182 222 40184 274
rect 40128 220 40184 222
rect 41188 274 41244 276
rect 41188 222 41190 274
rect 41190 222 41242 274
rect 41242 222 41244 274
rect 41188 220 41244 222
rect 1904 150 1960 152
rect 1904 98 1906 150
rect 1906 98 1958 150
rect 1958 98 1960 150
rect 1904 96 1960 98
rect 2036 150 2092 152
rect 2036 98 2038 150
rect 2038 98 2090 150
rect 2090 98 2092 150
rect 2036 96 2092 98
rect 3152 150 3208 152
rect 3152 98 3154 150
rect 3154 98 3206 150
rect 3206 98 3208 150
rect 3152 96 3208 98
rect 3284 150 3340 152
rect 3284 98 3286 150
rect 3286 98 3338 150
rect 3338 98 3340 150
rect 3284 96 3340 98
rect 4400 150 4456 152
rect 4400 98 4402 150
rect 4402 98 4454 150
rect 4454 98 4456 150
rect 4400 96 4456 98
rect 4532 150 4588 152
rect 4532 98 4534 150
rect 4534 98 4586 150
rect 4586 98 4588 150
rect 4532 96 4588 98
rect 5648 150 5704 152
rect 5648 98 5650 150
rect 5650 98 5702 150
rect 5702 98 5704 150
rect 5648 96 5704 98
rect 5780 150 5836 152
rect 5780 98 5782 150
rect 5782 98 5834 150
rect 5834 98 5836 150
rect 5780 96 5836 98
rect 6896 150 6952 152
rect 6896 98 6898 150
rect 6898 98 6950 150
rect 6950 98 6952 150
rect 6896 96 6952 98
rect 7028 150 7084 152
rect 7028 98 7030 150
rect 7030 98 7082 150
rect 7082 98 7084 150
rect 7028 96 7084 98
rect 8144 150 8200 152
rect 8144 98 8146 150
rect 8146 98 8198 150
rect 8198 98 8200 150
rect 8144 96 8200 98
rect 8276 150 8332 152
rect 8276 98 8278 150
rect 8278 98 8330 150
rect 8330 98 8332 150
rect 8276 96 8332 98
rect 9392 150 9448 152
rect 9392 98 9394 150
rect 9394 98 9446 150
rect 9446 98 9448 150
rect 9392 96 9448 98
rect 9524 150 9580 152
rect 9524 98 9526 150
rect 9526 98 9578 150
rect 9578 98 9580 150
rect 9524 96 9580 98
rect 10640 150 10696 152
rect 10640 98 10642 150
rect 10642 98 10694 150
rect 10694 98 10696 150
rect 10640 96 10696 98
rect 10772 150 10828 152
rect 10772 98 10774 150
rect 10774 98 10826 150
rect 10826 98 10828 150
rect 10772 96 10828 98
rect 11888 150 11944 152
rect 11888 98 11890 150
rect 11890 98 11942 150
rect 11942 98 11944 150
rect 11888 96 11944 98
rect 12020 150 12076 152
rect 12020 98 12022 150
rect 12022 98 12074 150
rect 12074 98 12076 150
rect 12020 96 12076 98
rect 13136 150 13192 152
rect 13136 98 13138 150
rect 13138 98 13190 150
rect 13190 98 13192 150
rect 13136 96 13192 98
rect 13268 150 13324 152
rect 13268 98 13270 150
rect 13270 98 13322 150
rect 13322 98 13324 150
rect 13268 96 13324 98
rect 14384 150 14440 152
rect 14384 98 14386 150
rect 14386 98 14438 150
rect 14438 98 14440 150
rect 14384 96 14440 98
rect 14516 150 14572 152
rect 14516 98 14518 150
rect 14518 98 14570 150
rect 14570 98 14572 150
rect 14516 96 14572 98
rect 15632 150 15688 152
rect 15632 98 15634 150
rect 15634 98 15686 150
rect 15686 98 15688 150
rect 15632 96 15688 98
rect 15764 150 15820 152
rect 15764 98 15766 150
rect 15766 98 15818 150
rect 15818 98 15820 150
rect 15764 96 15820 98
rect 16880 150 16936 152
rect 16880 98 16882 150
rect 16882 98 16934 150
rect 16934 98 16936 150
rect 16880 96 16936 98
rect 17012 150 17068 152
rect 17012 98 17014 150
rect 17014 98 17066 150
rect 17066 98 17068 150
rect 17012 96 17068 98
rect 18128 150 18184 152
rect 18128 98 18130 150
rect 18130 98 18182 150
rect 18182 98 18184 150
rect 18128 96 18184 98
rect 18260 150 18316 152
rect 18260 98 18262 150
rect 18262 98 18314 150
rect 18314 98 18316 150
rect 18260 96 18316 98
rect 19376 150 19432 152
rect 19376 98 19378 150
rect 19378 98 19430 150
rect 19430 98 19432 150
rect 19376 96 19432 98
rect 19508 150 19564 152
rect 19508 98 19510 150
rect 19510 98 19562 150
rect 19562 98 19564 150
rect 19508 96 19564 98
rect 20624 150 20680 152
rect 20624 98 20626 150
rect 20626 98 20678 150
rect 20678 98 20680 150
rect 20624 96 20680 98
rect 20756 150 20812 152
rect 20756 98 20758 150
rect 20758 98 20810 150
rect 20810 98 20812 150
rect 20756 96 20812 98
rect 21872 150 21928 152
rect 21872 98 21874 150
rect 21874 98 21926 150
rect 21926 98 21928 150
rect 21872 96 21928 98
rect 22004 150 22060 152
rect 22004 98 22006 150
rect 22006 98 22058 150
rect 22058 98 22060 150
rect 22004 96 22060 98
rect 23120 150 23176 152
rect 23120 98 23122 150
rect 23122 98 23174 150
rect 23174 98 23176 150
rect 23120 96 23176 98
rect 23252 150 23308 152
rect 23252 98 23254 150
rect 23254 98 23306 150
rect 23306 98 23308 150
rect 23252 96 23308 98
rect 24368 150 24424 152
rect 24368 98 24370 150
rect 24370 98 24422 150
rect 24422 98 24424 150
rect 24368 96 24424 98
rect 24500 150 24556 152
rect 24500 98 24502 150
rect 24502 98 24554 150
rect 24554 98 24556 150
rect 24500 96 24556 98
rect 25616 150 25672 152
rect 25616 98 25618 150
rect 25618 98 25670 150
rect 25670 98 25672 150
rect 25616 96 25672 98
rect 25748 150 25804 152
rect 25748 98 25750 150
rect 25750 98 25802 150
rect 25802 98 25804 150
rect 25748 96 25804 98
rect 26864 150 26920 152
rect 26864 98 26866 150
rect 26866 98 26918 150
rect 26918 98 26920 150
rect 26864 96 26920 98
rect 26996 150 27052 152
rect 26996 98 26998 150
rect 26998 98 27050 150
rect 27050 98 27052 150
rect 26996 96 27052 98
rect 28112 150 28168 152
rect 28112 98 28114 150
rect 28114 98 28166 150
rect 28166 98 28168 150
rect 28112 96 28168 98
rect 28244 150 28300 152
rect 28244 98 28246 150
rect 28246 98 28298 150
rect 28298 98 28300 150
rect 28244 96 28300 98
rect 29360 150 29416 152
rect 29360 98 29362 150
rect 29362 98 29414 150
rect 29414 98 29416 150
rect 29360 96 29416 98
rect 29492 150 29548 152
rect 29492 98 29494 150
rect 29494 98 29546 150
rect 29546 98 29548 150
rect 29492 96 29548 98
rect 30608 150 30664 152
rect 30608 98 30610 150
rect 30610 98 30662 150
rect 30662 98 30664 150
rect 30608 96 30664 98
rect 30740 150 30796 152
rect 30740 98 30742 150
rect 30742 98 30794 150
rect 30794 98 30796 150
rect 30740 96 30796 98
rect 31856 150 31912 152
rect 31856 98 31858 150
rect 31858 98 31910 150
rect 31910 98 31912 150
rect 31856 96 31912 98
rect 31988 150 32044 152
rect 31988 98 31990 150
rect 31990 98 32042 150
rect 32042 98 32044 150
rect 31988 96 32044 98
rect 33104 150 33160 152
rect 33104 98 33106 150
rect 33106 98 33158 150
rect 33158 98 33160 150
rect 33104 96 33160 98
rect 33236 150 33292 152
rect 33236 98 33238 150
rect 33238 98 33290 150
rect 33290 98 33292 150
rect 33236 96 33292 98
rect 34352 150 34408 152
rect 34352 98 34354 150
rect 34354 98 34406 150
rect 34406 98 34408 150
rect 34352 96 34408 98
rect 34484 150 34540 152
rect 34484 98 34486 150
rect 34486 98 34538 150
rect 34538 98 34540 150
rect 34484 96 34540 98
rect 35600 150 35656 152
rect 35600 98 35602 150
rect 35602 98 35654 150
rect 35654 98 35656 150
rect 35600 96 35656 98
rect 35732 150 35788 152
rect 35732 98 35734 150
rect 35734 98 35786 150
rect 35786 98 35788 150
rect 35732 96 35788 98
rect 36848 150 36904 152
rect 36848 98 36850 150
rect 36850 98 36902 150
rect 36902 98 36904 150
rect 36848 96 36904 98
rect 36980 150 37036 152
rect 36980 98 36982 150
rect 36982 98 37034 150
rect 37034 98 37036 150
rect 36980 96 37036 98
rect 38096 150 38152 152
rect 38096 98 38098 150
rect 38098 98 38150 150
rect 38150 98 38152 150
rect 38096 96 38152 98
rect 38228 150 38284 152
rect 38228 98 38230 150
rect 38230 98 38282 150
rect 38282 98 38284 150
rect 38228 96 38284 98
rect 39344 150 39400 152
rect 39344 98 39346 150
rect 39346 98 39398 150
rect 39398 98 39400 150
rect 39344 96 39400 98
rect 39476 150 39532 152
rect 39476 98 39478 150
rect 39478 98 39530 150
rect 39530 98 39532 150
rect 39476 96 39532 98
rect 40592 150 40648 152
rect 40592 98 40594 150
rect 40594 98 40646 150
rect 40646 98 40648 150
rect 40592 96 40648 98
rect 40724 150 40780 152
rect 40724 98 40726 150
rect 40726 98 40778 150
rect 40778 98 40780 150
rect 40724 96 40780 98
<< metal3 >>
rect 1949 1978 2047 2076
rect 3197 1978 3295 2076
rect 4445 1978 4543 2076
rect 5693 1978 5791 2076
rect 6941 1978 7039 2076
rect 8189 1978 8287 2076
rect 9437 1978 9535 2076
rect 10685 1978 10783 2076
rect 11933 1978 12031 2076
rect 13181 1978 13279 2076
rect 14429 1978 14527 2076
rect 15677 1978 15775 2076
rect 16925 1978 17023 2076
rect 18173 1978 18271 2076
rect 19421 1978 19519 2076
rect 20669 1978 20767 2076
rect 21917 1978 22015 2076
rect 23165 1978 23263 2076
rect 24413 1978 24511 2076
rect 25661 1978 25759 2076
rect 26909 1978 27007 2076
rect 28157 1978 28255 2076
rect 29405 1978 29503 2076
rect 30653 1978 30751 2076
rect 31901 1978 31999 2076
rect 33149 1978 33247 2076
rect 34397 1978 34495 2076
rect 35645 1978 35743 2076
rect 36893 1978 36991 2076
rect 38141 1978 38239 2076
rect 39389 1978 39487 2076
rect 40637 1978 40735 2076
rect 6021 1300 6087 1303
rect 11013 1300 11079 1303
rect 16005 1300 16071 1303
rect 20997 1300 21063 1303
rect 25989 1300 26055 1303
rect 30981 1300 31047 1303
rect 35973 1300 36039 1303
rect 40965 1300 41031 1303
rect 0 1298 41310 1300
rect 0 1242 6026 1298
rect 6082 1242 11018 1298
rect 11074 1242 16010 1298
rect 16066 1242 21002 1298
rect 21058 1242 25994 1298
rect 26050 1242 30986 1298
rect 31042 1242 35978 1298
rect 36034 1242 40970 1298
rect 41026 1242 41310 1298
rect 0 1240 41310 1242
rect 6021 1237 6087 1240
rect 11013 1237 11079 1240
rect 16005 1237 16071 1240
rect 20997 1237 21063 1240
rect 25989 1237 26055 1240
rect 30981 1237 31047 1240
rect 35973 1237 36039 1240
rect 40965 1237 41031 1240
rect 5397 1176 5463 1179
rect 10389 1176 10455 1179
rect 15381 1176 15447 1179
rect 20373 1176 20439 1179
rect 25365 1176 25431 1179
rect 30357 1176 30423 1179
rect 35349 1176 35415 1179
rect 40341 1176 40407 1179
rect 0 1174 41310 1176
rect 0 1118 5402 1174
rect 5458 1118 10394 1174
rect 10450 1118 15386 1174
rect 15442 1118 20378 1174
rect 20434 1118 25370 1174
rect 25426 1118 30362 1174
rect 30418 1118 35354 1174
rect 35410 1118 40346 1174
rect 40402 1118 41310 1174
rect 0 1116 41310 1118
rect 5397 1113 5463 1116
rect 10389 1113 10455 1116
rect 15381 1113 15447 1116
rect 20373 1113 20439 1116
rect 25365 1113 25431 1116
rect 30357 1113 30423 1116
rect 35349 1113 35415 1116
rect 40341 1113 40407 1116
rect 4773 1052 4839 1055
rect 9765 1052 9831 1055
rect 14757 1052 14823 1055
rect 19749 1052 19815 1055
rect 24741 1052 24807 1055
rect 29733 1052 29799 1055
rect 34725 1052 34791 1055
rect 39717 1052 39783 1055
rect 0 1050 41310 1052
rect 0 994 4778 1050
rect 4834 994 9770 1050
rect 9826 994 14762 1050
rect 14818 994 19754 1050
rect 19810 994 24746 1050
rect 24802 994 29738 1050
rect 29794 994 34730 1050
rect 34786 994 39722 1050
rect 39778 994 41310 1050
rect 0 992 41310 994
rect 4773 989 4839 992
rect 9765 989 9831 992
rect 14757 989 14823 992
rect 19749 989 19815 992
rect 24741 989 24807 992
rect 29733 989 29799 992
rect 34725 989 34791 992
rect 39717 989 39783 992
rect 4149 928 4215 931
rect 9141 928 9207 931
rect 14133 928 14199 931
rect 19125 928 19191 931
rect 24117 928 24183 931
rect 29109 928 29175 931
rect 34101 928 34167 931
rect 39093 928 39159 931
rect 0 926 41310 928
rect 0 870 4154 926
rect 4210 870 9146 926
rect 9202 870 14138 926
rect 14194 870 19130 926
rect 19186 870 24122 926
rect 24178 870 29114 926
rect 29170 870 34106 926
rect 34162 870 39098 926
rect 39154 870 41310 926
rect 0 868 41310 870
rect 4149 865 4215 868
rect 9141 865 9207 868
rect 14133 865 14199 868
rect 19125 865 19191 868
rect 24117 865 24183 868
rect 29109 865 29175 868
rect 34101 865 34167 868
rect 39093 865 39159 868
rect 3525 804 3591 807
rect 8517 804 8583 807
rect 13509 804 13575 807
rect 18501 804 18567 807
rect 23493 804 23559 807
rect 28485 804 28551 807
rect 33477 804 33543 807
rect 38469 804 38535 807
rect 0 802 41310 804
rect 0 746 3530 802
rect 3586 746 8522 802
rect 8578 746 13514 802
rect 13570 746 18506 802
rect 18562 746 23498 802
rect 23554 746 28490 802
rect 28546 746 33482 802
rect 33538 746 38474 802
rect 38530 746 41310 802
rect 0 744 41310 746
rect 3525 741 3591 744
rect 8517 741 8583 744
rect 13509 741 13575 744
rect 18501 741 18567 744
rect 23493 741 23559 744
rect 28485 741 28551 744
rect 33477 741 33543 744
rect 38469 741 38535 744
rect 2901 680 2967 683
rect 7893 680 7959 683
rect 12885 680 12951 683
rect 17877 680 17943 683
rect 22869 680 22935 683
rect 27861 680 27927 683
rect 32853 680 32919 683
rect 37845 680 37911 683
rect 0 678 41310 680
rect 0 622 2906 678
rect 2962 622 7898 678
rect 7954 622 12890 678
rect 12946 622 17882 678
rect 17938 622 22874 678
rect 22930 622 27866 678
rect 27922 622 32858 678
rect 32914 622 37850 678
rect 37906 622 41310 678
rect 0 620 41310 622
rect 2901 617 2967 620
rect 7893 617 7959 620
rect 12885 617 12951 620
rect 17877 617 17943 620
rect 22869 617 22935 620
rect 27861 617 27927 620
rect 32853 617 32919 620
rect 37845 617 37911 620
rect 2277 556 2343 559
rect 7269 556 7335 559
rect 12261 556 12327 559
rect 17253 556 17319 559
rect 22245 556 22311 559
rect 27237 556 27303 559
rect 32229 556 32295 559
rect 37221 556 37287 559
rect 0 554 41310 556
rect 0 498 2282 554
rect 2338 498 7274 554
rect 7330 498 12266 554
rect 12322 498 17258 554
rect 17314 498 22250 554
rect 22306 498 27242 554
rect 27298 498 32234 554
rect 32290 498 37226 554
rect 37282 498 41310 554
rect 0 496 41310 498
rect 2277 493 2343 496
rect 7269 493 7335 496
rect 12261 493 12327 496
rect 17253 493 17319 496
rect 22245 493 22311 496
rect 27237 493 27303 496
rect 32229 493 32295 496
rect 37221 493 37287 496
rect 1653 432 1719 435
rect 6645 432 6711 435
rect 11637 432 11703 435
rect 16629 432 16695 435
rect 21621 432 21687 435
rect 26613 432 26679 435
rect 31605 432 31671 435
rect 36597 432 36663 435
rect 0 430 41310 432
rect 0 374 1658 430
rect 1714 374 6650 430
rect 6706 374 11642 430
rect 11698 374 16634 430
rect 16690 374 21626 430
rect 21682 374 26618 430
rect 26674 374 31610 430
rect 31666 374 36602 430
rect 36658 374 41310 430
rect 0 372 41310 374
rect 1653 369 1719 372
rect 6645 369 6711 372
rect 11637 369 11703 372
rect 16629 369 16695 372
rect 21621 369 21687 372
rect 26613 369 26679 372
rect 31605 369 31671 372
rect 36597 369 36663 372
rect 1435 278 1501 281
rect 2495 278 2561 281
rect 2683 278 2749 281
rect 3743 278 3809 281
rect 3931 278 3997 281
rect 4991 278 5057 281
rect 5179 278 5245 281
rect 6239 278 6305 281
rect 1435 276 6305 278
rect 1435 220 1440 276
rect 1496 220 2500 276
rect 2556 220 2688 276
rect 2744 220 3748 276
rect 3804 220 3936 276
rect 3992 220 4996 276
rect 5052 220 5184 276
rect 5240 220 6244 276
rect 6300 220 6305 276
rect 1435 218 6305 220
rect 1435 215 1501 218
rect 2495 215 2561 218
rect 2683 215 2749 218
rect 3743 215 3809 218
rect 3931 215 3997 218
rect 4991 215 5057 218
rect 5179 215 5245 218
rect 6239 215 6305 218
rect 6427 278 6493 281
rect 7487 278 7553 281
rect 7675 278 7741 281
rect 8735 278 8801 281
rect 8923 278 8989 281
rect 9983 278 10049 281
rect 10171 278 10237 281
rect 11231 278 11297 281
rect 6427 276 11297 278
rect 6427 220 6432 276
rect 6488 220 7492 276
rect 7548 220 7680 276
rect 7736 220 8740 276
rect 8796 220 8928 276
rect 8984 220 9988 276
rect 10044 220 10176 276
rect 10232 220 11236 276
rect 11292 220 11297 276
rect 6427 218 11297 220
rect 6427 215 6493 218
rect 7487 215 7553 218
rect 7675 215 7741 218
rect 8735 215 8801 218
rect 8923 215 8989 218
rect 9983 215 10049 218
rect 10171 215 10237 218
rect 11231 215 11297 218
rect 11419 278 11485 281
rect 12479 278 12545 281
rect 12667 278 12733 281
rect 13727 278 13793 281
rect 13915 278 13981 281
rect 14975 278 15041 281
rect 15163 278 15229 281
rect 16223 278 16289 281
rect 11419 276 16289 278
rect 11419 220 11424 276
rect 11480 220 12484 276
rect 12540 220 12672 276
rect 12728 220 13732 276
rect 13788 220 13920 276
rect 13976 220 14980 276
rect 15036 220 15168 276
rect 15224 220 16228 276
rect 16284 220 16289 276
rect 11419 218 16289 220
rect 11419 215 11485 218
rect 12479 215 12545 218
rect 12667 215 12733 218
rect 13727 215 13793 218
rect 13915 215 13981 218
rect 14975 215 15041 218
rect 15163 215 15229 218
rect 16223 215 16289 218
rect 16411 278 16477 281
rect 17471 278 17537 281
rect 17659 278 17725 281
rect 18719 278 18785 281
rect 18907 278 18973 281
rect 19967 278 20033 281
rect 20155 278 20221 281
rect 21215 278 21281 281
rect 16411 276 21281 278
rect 16411 220 16416 276
rect 16472 220 17476 276
rect 17532 220 17664 276
rect 17720 220 18724 276
rect 18780 220 18912 276
rect 18968 220 19972 276
rect 20028 220 20160 276
rect 20216 220 21220 276
rect 21276 220 21281 276
rect 16411 218 21281 220
rect 16411 215 16477 218
rect 17471 215 17537 218
rect 17659 215 17725 218
rect 18719 215 18785 218
rect 18907 215 18973 218
rect 19967 215 20033 218
rect 20155 215 20221 218
rect 21215 215 21281 218
rect 21403 278 21469 281
rect 22463 278 22529 281
rect 22651 278 22717 281
rect 23711 278 23777 281
rect 23899 278 23965 281
rect 24959 278 25025 281
rect 25147 278 25213 281
rect 26207 278 26273 281
rect 21403 276 26273 278
rect 21403 220 21408 276
rect 21464 220 22468 276
rect 22524 220 22656 276
rect 22712 220 23716 276
rect 23772 220 23904 276
rect 23960 220 24964 276
rect 25020 220 25152 276
rect 25208 220 26212 276
rect 26268 220 26273 276
rect 21403 218 26273 220
rect 21403 215 21469 218
rect 22463 215 22529 218
rect 22651 215 22717 218
rect 23711 215 23777 218
rect 23899 215 23965 218
rect 24959 215 25025 218
rect 25147 215 25213 218
rect 26207 215 26273 218
rect 26395 278 26461 281
rect 27455 278 27521 281
rect 27643 278 27709 281
rect 28703 278 28769 281
rect 28891 278 28957 281
rect 29951 278 30017 281
rect 30139 278 30205 281
rect 31199 278 31265 281
rect 26395 276 31265 278
rect 26395 220 26400 276
rect 26456 220 27460 276
rect 27516 220 27648 276
rect 27704 220 28708 276
rect 28764 220 28896 276
rect 28952 220 29956 276
rect 30012 220 30144 276
rect 30200 220 31204 276
rect 31260 220 31265 276
rect 26395 218 31265 220
rect 26395 215 26461 218
rect 27455 215 27521 218
rect 27643 215 27709 218
rect 28703 215 28769 218
rect 28891 215 28957 218
rect 29951 215 30017 218
rect 30139 215 30205 218
rect 31199 215 31265 218
rect 31387 278 31453 281
rect 32447 278 32513 281
rect 32635 278 32701 281
rect 33695 278 33761 281
rect 33883 278 33949 281
rect 34943 278 35009 281
rect 35131 278 35197 281
rect 36191 278 36257 281
rect 31387 276 36257 278
rect 31387 220 31392 276
rect 31448 220 32452 276
rect 32508 220 32640 276
rect 32696 220 33700 276
rect 33756 220 33888 276
rect 33944 220 34948 276
rect 35004 220 35136 276
rect 35192 220 36196 276
rect 36252 220 36257 276
rect 31387 218 36257 220
rect 31387 215 31453 218
rect 32447 215 32513 218
rect 32635 215 32701 218
rect 33695 215 33761 218
rect 33883 215 33949 218
rect 34943 215 35009 218
rect 35131 215 35197 218
rect 36191 215 36257 218
rect 36379 278 36445 281
rect 37439 278 37505 281
rect 37627 278 37693 281
rect 38687 278 38753 281
rect 38875 278 38941 281
rect 39935 278 40001 281
rect 40123 278 40189 281
rect 41183 278 41249 281
rect 36379 276 41249 278
rect 36379 220 36384 276
rect 36440 220 37444 276
rect 37500 220 37632 276
rect 37688 220 38692 276
rect 38748 220 38880 276
rect 38936 220 39940 276
rect 39996 220 40128 276
rect 40184 220 41188 276
rect 41244 220 41249 276
rect 36379 218 41249 220
rect 36379 215 36445 218
rect 37439 215 37505 218
rect 37627 215 37693 218
rect 38687 215 38753 218
rect 38875 215 38941 218
rect 39935 215 40001 218
rect 40123 215 40189 218
rect 41183 215 41249 218
rect 1899 154 1965 157
rect 2031 154 2097 157
rect 3147 154 3213 157
rect 3279 154 3345 157
rect 4395 154 4461 157
rect 4527 154 4593 157
rect 5643 154 5709 157
rect 5775 154 5841 157
rect 1899 152 5841 154
rect 1899 96 1904 152
rect 1960 96 2036 152
rect 2092 96 3152 152
rect 3208 96 3284 152
rect 3340 96 4400 152
rect 4456 96 4532 152
rect 4588 96 5648 152
rect 5704 96 5780 152
rect 5836 96 5841 152
rect 1899 94 5841 96
rect 1899 91 1965 94
rect 2031 91 2097 94
rect 3147 91 3213 94
rect 3279 91 3345 94
rect 4395 91 4461 94
rect 4527 91 4593 94
rect 5643 91 5709 94
rect 5775 91 5841 94
rect 6891 154 6957 157
rect 7023 154 7089 157
rect 8139 154 8205 157
rect 8271 154 8337 157
rect 9387 154 9453 157
rect 9519 154 9585 157
rect 10635 154 10701 157
rect 10767 154 10833 157
rect 6891 152 10833 154
rect 6891 96 6896 152
rect 6952 96 7028 152
rect 7084 96 8144 152
rect 8200 96 8276 152
rect 8332 96 9392 152
rect 9448 96 9524 152
rect 9580 96 10640 152
rect 10696 96 10772 152
rect 10828 96 10833 152
rect 6891 94 10833 96
rect 6891 91 6957 94
rect 7023 91 7089 94
rect 8139 91 8205 94
rect 8271 91 8337 94
rect 9387 91 9453 94
rect 9519 91 9585 94
rect 10635 91 10701 94
rect 10767 91 10833 94
rect 11883 154 11949 157
rect 12015 154 12081 157
rect 13131 154 13197 157
rect 13263 154 13329 157
rect 14379 154 14445 157
rect 14511 154 14577 157
rect 15627 154 15693 157
rect 15759 154 15825 157
rect 11883 152 15825 154
rect 11883 96 11888 152
rect 11944 96 12020 152
rect 12076 96 13136 152
rect 13192 96 13268 152
rect 13324 96 14384 152
rect 14440 96 14516 152
rect 14572 96 15632 152
rect 15688 96 15764 152
rect 15820 96 15825 152
rect 11883 94 15825 96
rect 11883 91 11949 94
rect 12015 91 12081 94
rect 13131 91 13197 94
rect 13263 91 13329 94
rect 14379 91 14445 94
rect 14511 91 14577 94
rect 15627 91 15693 94
rect 15759 91 15825 94
rect 16875 154 16941 157
rect 17007 154 17073 157
rect 18123 154 18189 157
rect 18255 154 18321 157
rect 19371 154 19437 157
rect 19503 154 19569 157
rect 20619 154 20685 157
rect 20751 154 20817 157
rect 16875 152 20817 154
rect 16875 96 16880 152
rect 16936 96 17012 152
rect 17068 96 18128 152
rect 18184 96 18260 152
rect 18316 96 19376 152
rect 19432 96 19508 152
rect 19564 96 20624 152
rect 20680 96 20756 152
rect 20812 96 20817 152
rect 16875 94 20817 96
rect 16875 91 16941 94
rect 17007 91 17073 94
rect 18123 91 18189 94
rect 18255 91 18321 94
rect 19371 91 19437 94
rect 19503 91 19569 94
rect 20619 91 20685 94
rect 20751 91 20817 94
rect 21867 154 21933 157
rect 21999 154 22065 157
rect 23115 154 23181 157
rect 23247 154 23313 157
rect 24363 154 24429 157
rect 24495 154 24561 157
rect 25611 154 25677 157
rect 25743 154 25809 157
rect 21867 152 25809 154
rect 21867 96 21872 152
rect 21928 96 22004 152
rect 22060 96 23120 152
rect 23176 96 23252 152
rect 23308 96 24368 152
rect 24424 96 24500 152
rect 24556 96 25616 152
rect 25672 96 25748 152
rect 25804 96 25809 152
rect 21867 94 25809 96
rect 21867 91 21933 94
rect 21999 91 22065 94
rect 23115 91 23181 94
rect 23247 91 23313 94
rect 24363 91 24429 94
rect 24495 91 24561 94
rect 25611 91 25677 94
rect 25743 91 25809 94
rect 26859 154 26925 157
rect 26991 154 27057 157
rect 28107 154 28173 157
rect 28239 154 28305 157
rect 29355 154 29421 157
rect 29487 154 29553 157
rect 30603 154 30669 157
rect 30735 154 30801 157
rect 26859 152 30801 154
rect 26859 96 26864 152
rect 26920 96 26996 152
rect 27052 96 28112 152
rect 28168 96 28244 152
rect 28300 96 29360 152
rect 29416 96 29492 152
rect 29548 96 30608 152
rect 30664 96 30740 152
rect 30796 96 30801 152
rect 26859 94 30801 96
rect 26859 91 26925 94
rect 26991 91 27057 94
rect 28107 91 28173 94
rect 28239 91 28305 94
rect 29355 91 29421 94
rect 29487 91 29553 94
rect 30603 91 30669 94
rect 30735 91 30801 94
rect 31851 154 31917 157
rect 31983 154 32049 157
rect 33099 154 33165 157
rect 33231 154 33297 157
rect 34347 154 34413 157
rect 34479 154 34545 157
rect 35595 154 35661 157
rect 35727 154 35793 157
rect 31851 152 35793 154
rect 31851 96 31856 152
rect 31912 96 31988 152
rect 32044 96 33104 152
rect 33160 96 33236 152
rect 33292 96 34352 152
rect 34408 96 34484 152
rect 34540 96 35600 152
rect 35656 96 35732 152
rect 35788 96 35793 152
rect 31851 94 35793 96
rect 31851 91 31917 94
rect 31983 91 32049 94
rect 33099 91 33165 94
rect 33231 91 33297 94
rect 34347 91 34413 94
rect 34479 91 34545 94
rect 35595 91 35661 94
rect 35727 91 35793 94
rect 36843 154 36909 157
rect 36975 154 37041 157
rect 38091 154 38157 157
rect 38223 154 38289 157
rect 39339 154 39405 157
rect 39471 154 39537 157
rect 40587 154 40653 157
rect 40719 154 40785 157
rect 36843 152 40785 154
rect 36843 96 36848 152
rect 36904 96 36980 152
rect 37036 96 38096 152
rect 38152 96 38228 152
rect 38284 96 39344 152
rect 39400 96 39476 152
rect 39532 96 40592 152
rect 40648 96 40724 152
rect 40780 96 40785 152
rect 36843 94 40785 96
rect 36843 91 36909 94
rect 36975 91 37041 94
rect 38091 91 38157 94
rect 38223 91 38289 94
rect 39339 91 39405 94
rect 39471 91 39537 94
rect 40587 91 40653 94
rect 40719 91 40785 94
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_0
timestamp 1723858470
transform -1 0 11358 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_1
timestamp 1723858470
transform 1 0 10110 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_2
timestamp 1723858470
transform -1 0 10110 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_3
timestamp 1723858470
transform 1 0 8862 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_4
timestamp 1723858470
transform -1 0 8862 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_5
timestamp 1723858470
transform 1 0 7614 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_6
timestamp 1723858470
transform -1 0 7614 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_7
timestamp 1723858470
transform 1 0 6366 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_8
timestamp 1723858470
transform -1 0 6366 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_9
timestamp 1723858470
transform 1 0 5118 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_10
timestamp 1723858470
transform -1 0 5118 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_11
timestamp 1723858470
transform 1 0 3870 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_12
timestamp 1723858470
transform -1 0 3870 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_13
timestamp 1723858470
transform 1 0 2622 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_14
timestamp 1723858470
transform -1 0 2622 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_15
timestamp 1723858470
transform 1 0 1374 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_16
timestamp 1723858470
transform -1 0 21342 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_17
timestamp 1723858470
transform 1 0 20094 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_18
timestamp 1723858470
transform -1 0 20094 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_19
timestamp 1723858470
transform 1 0 18846 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_20
timestamp 1723858470
transform -1 0 18846 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_21
timestamp 1723858470
transform 1 0 17598 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_22
timestamp 1723858470
transform -1 0 17598 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_23
timestamp 1723858470
transform 1 0 16350 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_24
timestamp 1723858470
transform -1 0 16350 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_25
timestamp 1723858470
transform 1 0 15102 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_26
timestamp 1723858470
transform -1 0 15102 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_27
timestamp 1723858470
transform 1 0 13854 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_28
timestamp 1723858470
transform -1 0 13854 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_29
timestamp 1723858470
transform 1 0 12606 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_30
timestamp 1723858470
transform -1 0 12606 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_31
timestamp 1723858470
transform 1 0 11358 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_32
timestamp 1723858470
transform -1 0 31326 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_33
timestamp 1723858470
transform 1 0 30078 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_34
timestamp 1723858470
transform -1 0 30078 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_35
timestamp 1723858470
transform 1 0 28830 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_36
timestamp 1723858470
transform -1 0 28830 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_37
timestamp 1723858470
transform 1 0 27582 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_38
timestamp 1723858470
transform -1 0 27582 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_39
timestamp 1723858470
transform 1 0 26334 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_40
timestamp 1723858470
transform -1 0 26334 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_41
timestamp 1723858470
transform 1 0 25086 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_42
timestamp 1723858470
transform -1 0 25086 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_43
timestamp 1723858470
transform 1 0 23838 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_44
timestamp 1723858470
transform -1 0 23838 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_45
timestamp 1723858470
transform 1 0 22590 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_46
timestamp 1723858470
transform -1 0 22590 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_47
timestamp 1723858470
transform 1 0 21342 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_48
timestamp 1723858470
transform -1 0 41310 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_49
timestamp 1723858470
transform 1 0 40062 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_50
timestamp 1723858470
transform -1 0 40062 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_51
timestamp 1723858470
transform 1 0 38814 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_52
timestamp 1723858470
transform -1 0 38814 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_53
timestamp 1723858470
transform 1 0 37566 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_54
timestamp 1723858470
transform -1 0 37566 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_55
timestamp 1723858470
transform 1 0 36318 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_56
timestamp 1723858470
transform -1 0 36318 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_57
timestamp 1723858470
transform 1 0 35070 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_58
timestamp 1723858470
transform -1 0 35070 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_59
timestamp 1723858470
transform 1 0 33822 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_60
timestamp 1723858470
transform -1 0 33822 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_61
timestamp 1723858470
transform 1 0 32574 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_62
timestamp 1723858470
transform -1 0 32574 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_63
timestamp 1723858470
transform 1 0 31326 0 1 1364
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_0
timestamp 1723858470
transform 1 0 11013 0 1 1237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_1
timestamp 1723858470
transform 1 0 10389 0 1 1113
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_2
timestamp 1723858470
transform 1 0 9765 0 1 989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_3
timestamp 1723858470
transform 1 0 9141 0 1 865
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_4
timestamp 1723858470
transform 1 0 8517 0 1 741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_5
timestamp 1723858470
transform 1 0 7893 0 1 617
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_6
timestamp 1723858470
transform 1 0 7269 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_7
timestamp 1723858470
transform 1 0 6645 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_8
timestamp 1723858470
transform 1 0 6021 0 1 1237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_9
timestamp 1723858470
transform 1 0 5397 0 1 1113
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_10
timestamp 1723858470
transform 1 0 4773 0 1 989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_11
timestamp 1723858470
transform 1 0 4149 0 1 865
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_12
timestamp 1723858470
transform 1 0 3525 0 1 741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_13
timestamp 1723858470
transform 1 0 2901 0 1 617
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_14
timestamp 1723858470
transform 1 0 2277 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_15
timestamp 1723858470
transform 1 0 1653 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_16
timestamp 1723858470
transform 1 0 20997 0 1 1237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_17
timestamp 1723858470
transform 1 0 20373 0 1 1113
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_18
timestamp 1723858470
transform 1 0 19749 0 1 989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_19
timestamp 1723858470
transform 1 0 19125 0 1 865
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_20
timestamp 1723858470
transform 1 0 18501 0 1 741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_21
timestamp 1723858470
transform 1 0 17877 0 1 617
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_22
timestamp 1723858470
transform 1 0 17253 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_23
timestamp 1723858470
transform 1 0 16629 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_24
timestamp 1723858470
transform 1 0 13509 0 1 741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_25
timestamp 1723858470
transform 1 0 12885 0 1 617
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_26
timestamp 1723858470
transform 1 0 12261 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_27
timestamp 1723858470
transform 1 0 11637 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_28
timestamp 1723858470
transform 1 0 16005 0 1 1237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_29
timestamp 1723858470
transform 1 0 15381 0 1 1113
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_30
timestamp 1723858470
transform 1 0 14757 0 1 989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_31
timestamp 1723858470
transform 1 0 14133 0 1 865
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_32
timestamp 1723858470
transform 1 0 28485 0 1 741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_33
timestamp 1723858470
transform 1 0 27861 0 1 617
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_34
timestamp 1723858470
transform 1 0 27237 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_35
timestamp 1723858470
transform 1 0 26613 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_36
timestamp 1723858470
transform 1 0 30981 0 1 1237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_37
timestamp 1723858470
transform 1 0 30357 0 1 1113
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_38
timestamp 1723858470
transform 1 0 29733 0 1 989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_39
timestamp 1723858470
transform 1 0 29109 0 1 865
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_40
timestamp 1723858470
transform 1 0 25989 0 1 1237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_41
timestamp 1723858470
transform 1 0 25365 0 1 1113
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_42
timestamp 1723858470
transform 1 0 24741 0 1 989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_43
timestamp 1723858470
transform 1 0 24117 0 1 865
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_44
timestamp 1723858470
transform 1 0 23493 0 1 741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_45
timestamp 1723858470
transform 1 0 22869 0 1 617
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_46
timestamp 1723858470
transform 1 0 22245 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_47
timestamp 1723858470
transform 1 0 21621 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_48
timestamp 1723858470
transform 1 0 40965 0 1 1237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_49
timestamp 1723858470
transform 1 0 40341 0 1 1113
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_50
timestamp 1723858470
transform 1 0 39717 0 1 989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_51
timestamp 1723858470
transform 1 0 39093 0 1 865
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_52
timestamp 1723858470
transform 1 0 38469 0 1 741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_53
timestamp 1723858470
transform 1 0 37845 0 1 617
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_54
timestamp 1723858470
transform 1 0 37221 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_55
timestamp 1723858470
transform 1 0 36597 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_56
timestamp 1723858470
transform 1 0 35973 0 1 1237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_57
timestamp 1723858470
transform 1 0 35349 0 1 1113
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_58
timestamp 1723858470
transform 1 0 34725 0 1 989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_59
timestamp 1723858470
transform 1 0 34101 0 1 865
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_60
timestamp 1723858470
transform 1 0 33477 0 1 741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_61
timestamp 1723858470
transform 1 0 32853 0 1 617
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_62
timestamp 1723858470
transform 1 0 32229 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_24_63
timestamp 1723858470
transform 1 0 31605 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_0
timestamp 1723858470
transform 1 0 11017 0 1 1237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_1
timestamp 1723858470
transform 1 0 10393 0 1 1113
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_2
timestamp 1723858470
transform 1 0 9769 0 1 989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_3
timestamp 1723858470
transform 1 0 9145 0 1 865
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_4
timestamp 1723858470
transform 1 0 8521 0 1 741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_5
timestamp 1723858470
transform 1 0 7897 0 1 617
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_6
timestamp 1723858470
transform 1 0 7273 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_7
timestamp 1723858470
transform 1 0 6649 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_8
timestamp 1723858470
transform 1 0 6025 0 1 1237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_9
timestamp 1723858470
transform 1 0 5401 0 1 1113
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_10
timestamp 1723858470
transform 1 0 4777 0 1 989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_11
timestamp 1723858470
transform 1 0 4153 0 1 865
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_12
timestamp 1723858470
transform 1 0 3529 0 1 741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_13
timestamp 1723858470
transform 1 0 2905 0 1 617
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_14
timestamp 1723858470
transform 1 0 2281 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_15
timestamp 1723858470
transform 1 0 1657 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_16
timestamp 1723858470
transform 1 0 21001 0 1 1237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_17
timestamp 1723858470
transform 1 0 20377 0 1 1113
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_18
timestamp 1723858470
transform 1 0 19753 0 1 989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_19
timestamp 1723858470
transform 1 0 19129 0 1 865
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_20
timestamp 1723858470
transform 1 0 18505 0 1 741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_21
timestamp 1723858470
transform 1 0 17881 0 1 617
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_22
timestamp 1723858470
transform 1 0 17257 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_23
timestamp 1723858470
transform 1 0 16633 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_24
timestamp 1723858470
transform 1 0 13513 0 1 741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_25
timestamp 1723858470
transform 1 0 12889 0 1 617
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_26
timestamp 1723858470
transform 1 0 12265 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_27
timestamp 1723858470
transform 1 0 11641 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_28
timestamp 1723858470
transform 1 0 16009 0 1 1237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_29
timestamp 1723858470
transform 1 0 15385 0 1 1113
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_30
timestamp 1723858470
transform 1 0 14761 0 1 989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_31
timestamp 1723858470
transform 1 0 14137 0 1 865
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_32
timestamp 1723858470
transform 1 0 28489 0 1 741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_33
timestamp 1723858470
transform 1 0 27865 0 1 617
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_34
timestamp 1723858470
transform 1 0 27241 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_35
timestamp 1723858470
transform 1 0 26617 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_36
timestamp 1723858470
transform 1 0 30985 0 1 1237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_37
timestamp 1723858470
transform 1 0 30361 0 1 1113
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_38
timestamp 1723858470
transform 1 0 29737 0 1 989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_39
timestamp 1723858470
transform 1 0 29113 0 1 865
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_40
timestamp 1723858470
transform 1 0 25993 0 1 1237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_41
timestamp 1723858470
transform 1 0 25369 0 1 1113
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_42
timestamp 1723858470
transform 1 0 24745 0 1 989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_43
timestamp 1723858470
transform 1 0 24121 0 1 865
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_44
timestamp 1723858470
transform 1 0 23497 0 1 741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_45
timestamp 1723858470
transform 1 0 22873 0 1 617
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_46
timestamp 1723858470
transform 1 0 22249 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_47
timestamp 1723858470
transform 1 0 21625 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_48
timestamp 1723858470
transform 1 0 40969 0 1 1237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_49
timestamp 1723858470
transform 1 0 40345 0 1 1113
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_50
timestamp 1723858470
transform 1 0 39721 0 1 989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_51
timestamp 1723858470
transform 1 0 39097 0 1 865
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_52
timestamp 1723858470
transform 1 0 38473 0 1 741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_53
timestamp 1723858470
transform 1 0 37849 0 1 617
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_54
timestamp 1723858470
transform 1 0 37225 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_55
timestamp 1723858470
transform 1 0 36601 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_56
timestamp 1723858470
transform 1 0 35977 0 1 1237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_57
timestamp 1723858470
transform 1 0 35353 0 1 1113
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_58
timestamp 1723858470
transform 1 0 34729 0 1 989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_59
timestamp 1723858470
transform 1 0 34105 0 1 865
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_60
timestamp 1723858470
transform 1 0 33481 0 1 741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_61
timestamp 1723858470
transform 1 0 32857 0 1 617
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_62
timestamp 1723858470
transform 1 0 32233 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_25_63
timestamp 1723858470
transform 1 0 31609 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_0
timestamp 1723858470
transform 1 0 11014 0 1 1238
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_1
timestamp 1723858470
transform 1 0 10390 0 1 1114
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_2
timestamp 1723858470
transform 1 0 9766 0 1 990
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_3
timestamp 1723858470
transform 1 0 9142 0 1 866
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_4
timestamp 1723858470
transform 1 0 8518 0 1 742
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_5
timestamp 1723858470
transform 1 0 7894 0 1 618
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_6
timestamp 1723858470
transform 1 0 7270 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_7
timestamp 1723858470
transform 1 0 6646 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_8
timestamp 1723858470
transform 1 0 8272 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_9
timestamp 1723858470
transform 1 0 8736 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_10
timestamp 1723858470
transform 1 0 8140 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_11
timestamp 1723858470
transform 1 0 7676 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_12
timestamp 1723858470
transform 1 0 7024 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_13
timestamp 1723858470
transform 1 0 7488 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_14
timestamp 1723858470
transform 1 0 6892 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_15
timestamp 1723858470
transform 1 0 6428 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_16
timestamp 1723858470
transform 1 0 10768 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_17
timestamp 1723858470
transform 1 0 11232 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_18
timestamp 1723858470
transform 1 0 10636 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_19
timestamp 1723858470
transform 1 0 10172 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_20
timestamp 1723858470
transform 1 0 9520 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_21
timestamp 1723858470
transform 1 0 9984 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_22
timestamp 1723858470
transform 1 0 9388 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_23
timestamp 1723858470
transform 1 0 8924 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_24
timestamp 1723858470
transform 1 0 6022 0 1 1238
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_25
timestamp 1723858470
transform 1 0 5398 0 1 1114
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_26
timestamp 1723858470
transform 1 0 4774 0 1 990
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_27
timestamp 1723858470
transform 1 0 4150 0 1 866
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_28
timestamp 1723858470
transform 1 0 3526 0 1 742
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_29
timestamp 1723858470
transform 1 0 2902 0 1 618
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_30
timestamp 1723858470
transform 1 0 2278 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_31
timestamp 1723858470
transform 1 0 1654 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_32
timestamp 1723858470
transform 1 0 3280 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_33
timestamp 1723858470
transform 1 0 3744 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_34
timestamp 1723858470
transform 1 0 3148 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_35
timestamp 1723858470
transform 1 0 2684 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_36
timestamp 1723858470
transform 1 0 2032 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_37
timestamp 1723858470
transform 1 0 2496 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_38
timestamp 1723858470
transform 1 0 1900 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_39
timestamp 1723858470
transform 1 0 1436 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_40
timestamp 1723858470
transform 1 0 5776 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_41
timestamp 1723858470
transform 1 0 6240 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_42
timestamp 1723858470
transform 1 0 5644 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_43
timestamp 1723858470
transform 1 0 5180 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_44
timestamp 1723858470
transform 1 0 4528 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_45
timestamp 1723858470
transform 1 0 4992 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_46
timestamp 1723858470
transform 1 0 4396 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_47
timestamp 1723858470
transform 1 0 3932 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_48
timestamp 1723858470
transform 1 0 18256 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_49
timestamp 1723858470
transform 1 0 18720 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_50
timestamp 1723858470
transform 1 0 18124 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_51
timestamp 1723858470
transform 1 0 17660 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_52
timestamp 1723858470
transform 1 0 17008 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_53
timestamp 1723858470
transform 1 0 17472 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_54
timestamp 1723858470
transform 1 0 16876 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_55
timestamp 1723858470
transform 1 0 16412 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_56
timestamp 1723858470
transform 1 0 20998 0 1 1238
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_57
timestamp 1723858470
transform 1 0 20374 0 1 1114
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_58
timestamp 1723858470
transform 1 0 19750 0 1 990
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_59
timestamp 1723858470
transform 1 0 19126 0 1 866
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_60
timestamp 1723858470
transform 1 0 18502 0 1 742
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_61
timestamp 1723858470
transform 1 0 17878 0 1 618
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_62
timestamp 1723858470
transform 1 0 17254 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_63
timestamp 1723858470
transform 1 0 16630 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_64
timestamp 1723858470
transform 1 0 20752 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_65
timestamp 1723858470
transform 1 0 21216 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_66
timestamp 1723858470
transform 1 0 20620 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_67
timestamp 1723858470
transform 1 0 20156 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_68
timestamp 1723858470
transform 1 0 19504 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_69
timestamp 1723858470
transform 1 0 19968 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_70
timestamp 1723858470
transform 1 0 19372 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_71
timestamp 1723858470
transform 1 0 18908 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_72
timestamp 1723858470
transform 1 0 13510 0 1 742
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_73
timestamp 1723858470
transform 1 0 12886 0 1 618
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_74
timestamp 1723858470
transform 1 0 12262 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_75
timestamp 1723858470
transform 1 0 11638 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_76
timestamp 1723858470
transform 1 0 15760 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_77
timestamp 1723858470
transform 1 0 16224 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_78
timestamp 1723858470
transform 1 0 15628 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_79
timestamp 1723858470
transform 1 0 15164 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_80
timestamp 1723858470
transform 1 0 14512 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_81
timestamp 1723858470
transform 1 0 14976 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_82
timestamp 1723858470
transform 1 0 14380 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_83
timestamp 1723858470
transform 1 0 13916 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_84
timestamp 1723858470
transform 1 0 13264 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_85
timestamp 1723858470
transform 1 0 13728 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_86
timestamp 1723858470
transform 1 0 13132 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_87
timestamp 1723858470
transform 1 0 12668 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_88
timestamp 1723858470
transform 1 0 12016 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_89
timestamp 1723858470
transform 1 0 12480 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_90
timestamp 1723858470
transform 1 0 11884 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_91
timestamp 1723858470
transform 1 0 11420 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_92
timestamp 1723858470
transform 1 0 16006 0 1 1238
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_93
timestamp 1723858470
transform 1 0 15382 0 1 1114
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_94
timestamp 1723858470
transform 1 0 14758 0 1 990
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_95
timestamp 1723858470
transform 1 0 14134 0 1 866
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_96
timestamp 1723858470
transform 1 0 30736 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_97
timestamp 1723858470
transform 1 0 31200 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_98
timestamp 1723858470
transform 1 0 30604 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_99
timestamp 1723858470
transform 1 0 30140 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_100
timestamp 1723858470
transform 1 0 29488 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_101
timestamp 1723858470
transform 1 0 29952 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_102
timestamp 1723858470
transform 1 0 29356 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_103
timestamp 1723858470
transform 1 0 28892 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_104
timestamp 1723858470
transform 1 0 28240 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_105
timestamp 1723858470
transform 1 0 28704 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_106
timestamp 1723858470
transform 1 0 28108 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_107
timestamp 1723858470
transform 1 0 27644 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_108
timestamp 1723858470
transform 1 0 26992 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_109
timestamp 1723858470
transform 1 0 27456 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_110
timestamp 1723858470
transform 1 0 26860 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_111
timestamp 1723858470
transform 1 0 26396 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_112
timestamp 1723858470
transform 1 0 28486 0 1 742
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_113
timestamp 1723858470
transform 1 0 27862 0 1 618
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_114
timestamp 1723858470
transform 1 0 27238 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_115
timestamp 1723858470
transform 1 0 26614 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_116
timestamp 1723858470
transform 1 0 30982 0 1 1238
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_117
timestamp 1723858470
transform 1 0 30358 0 1 1114
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_118
timestamp 1723858470
transform 1 0 29734 0 1 990
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_119
timestamp 1723858470
transform 1 0 29110 0 1 866
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_120
timestamp 1723858470
transform 1 0 25990 0 1 1238
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_121
timestamp 1723858470
transform 1 0 25366 0 1 1114
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_122
timestamp 1723858470
transform 1 0 24742 0 1 990
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_123
timestamp 1723858470
transform 1 0 24118 0 1 866
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_124
timestamp 1723858470
transform 1 0 23494 0 1 742
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_125
timestamp 1723858470
transform 1 0 22870 0 1 618
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_126
timestamp 1723858470
transform 1 0 22246 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_127
timestamp 1723858470
transform 1 0 21622 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_128
timestamp 1723858470
transform 1 0 23248 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_129
timestamp 1723858470
transform 1 0 23712 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_130
timestamp 1723858470
transform 1 0 23116 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_131
timestamp 1723858470
transform 1 0 22652 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_132
timestamp 1723858470
transform 1 0 22000 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_133
timestamp 1723858470
transform 1 0 22464 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_134
timestamp 1723858470
transform 1 0 21868 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_135
timestamp 1723858470
transform 1 0 21404 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_136
timestamp 1723858470
transform 1 0 25744 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_137
timestamp 1723858470
transform 1 0 26208 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_138
timestamp 1723858470
transform 1 0 25612 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_139
timestamp 1723858470
transform 1 0 25148 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_140
timestamp 1723858470
transform 1 0 24496 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_141
timestamp 1723858470
transform 1 0 24960 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_142
timestamp 1723858470
transform 1 0 24364 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_143
timestamp 1723858470
transform 1 0 23900 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_144
timestamp 1723858470
transform 1 0 40720 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_145
timestamp 1723858470
transform 1 0 41184 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_146
timestamp 1723858470
transform 1 0 40588 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_147
timestamp 1723858470
transform 1 0 40124 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_148
timestamp 1723858470
transform 1 0 39472 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_149
timestamp 1723858470
transform 1 0 39936 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_150
timestamp 1723858470
transform 1 0 39340 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_151
timestamp 1723858470
transform 1 0 38876 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_152
timestamp 1723858470
transform 1 0 38224 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_153
timestamp 1723858470
transform 1 0 38688 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_154
timestamp 1723858470
transform 1 0 38092 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_155
timestamp 1723858470
transform 1 0 37628 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_156
timestamp 1723858470
transform 1 0 36976 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_157
timestamp 1723858470
transform 1 0 37440 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_158
timestamp 1723858470
transform 1 0 36844 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_159
timestamp 1723858470
transform 1 0 36380 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_160
timestamp 1723858470
transform 1 0 40966 0 1 1238
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_161
timestamp 1723858470
transform 1 0 40342 0 1 1114
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_162
timestamp 1723858470
transform 1 0 39718 0 1 990
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_163
timestamp 1723858470
transform 1 0 39094 0 1 866
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_164
timestamp 1723858470
transform 1 0 38470 0 1 742
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_165
timestamp 1723858470
transform 1 0 37846 0 1 618
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_166
timestamp 1723858470
transform 1 0 37222 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_167
timestamp 1723858470
transform 1 0 36598 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_168
timestamp 1723858470
transform 1 0 35728 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_169
timestamp 1723858470
transform 1 0 36192 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_170
timestamp 1723858470
transform 1 0 35596 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_171
timestamp 1723858470
transform 1 0 35132 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_172
timestamp 1723858470
transform 1 0 34480 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_173
timestamp 1723858470
transform 1 0 34944 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_174
timestamp 1723858470
transform 1 0 34348 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_175
timestamp 1723858470
transform 1 0 33884 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_176
timestamp 1723858470
transform 1 0 33232 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_177
timestamp 1723858470
transform 1 0 33696 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_178
timestamp 1723858470
transform 1 0 33100 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_179
timestamp 1723858470
transform 1 0 32636 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_180
timestamp 1723858470
transform 1 0 31984 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_181
timestamp 1723858470
transform 1 0 32448 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_182
timestamp 1723858470
transform 1 0 31852 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_183
timestamp 1723858470
transform 1 0 31388 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_184
timestamp 1723858470
transform 1 0 35974 0 1 1238
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_185
timestamp 1723858470
transform 1 0 35350 0 1 1114
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_186
timestamp 1723858470
transform 1 0 34726 0 1 990
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_187
timestamp 1723858470
transform 1 0 34102 0 1 866
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_188
timestamp 1723858470
transform 1 0 33478 0 1 742
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_189
timestamp 1723858470
transform 1 0 32854 0 1 618
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_190
timestamp 1723858470
transform 1 0 32230 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_26_191
timestamp 1723858470
transform 1 0 31606 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_0
timestamp 1723858470
transform 1 0 11013 0 1 1233
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_1
timestamp 1723858470
transform 1 0 10389 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_2
timestamp 1723858470
transform 1 0 9765 0 1 985
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_3
timestamp 1723858470
transform 1 0 9141 0 1 861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_4
timestamp 1723858470
transform 1 0 8517 0 1 737
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_5
timestamp 1723858470
transform 1 0 7893 0 1 613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_6
timestamp 1723858470
transform 1 0 7269 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_7
timestamp 1723858470
transform 1 0 6645 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_8
timestamp 1723858470
transform 1 0 8271 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_9
timestamp 1723858470
transform 1 0 8735 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_10
timestamp 1723858470
transform 1 0 8139 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_11
timestamp 1723858470
transform 1 0 7675 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_12
timestamp 1723858470
transform 1 0 7023 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_13
timestamp 1723858470
transform 1 0 7487 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_14
timestamp 1723858470
transform 1 0 6891 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_15
timestamp 1723858470
transform 1 0 6427 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_16
timestamp 1723858470
transform 1 0 10767 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_17
timestamp 1723858470
transform 1 0 11231 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_18
timestamp 1723858470
transform 1 0 10635 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_19
timestamp 1723858470
transform 1 0 10171 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_20
timestamp 1723858470
transform 1 0 9519 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_21
timestamp 1723858470
transform 1 0 9983 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_22
timestamp 1723858470
transform 1 0 9387 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_23
timestamp 1723858470
transform 1 0 8923 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_24
timestamp 1723858470
transform 1 0 6021 0 1 1233
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_25
timestamp 1723858470
transform 1 0 5397 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_26
timestamp 1723858470
transform 1 0 4773 0 1 985
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_27
timestamp 1723858470
transform 1 0 4149 0 1 861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_28
timestamp 1723858470
transform 1 0 3525 0 1 737
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_29
timestamp 1723858470
transform 1 0 2901 0 1 613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_30
timestamp 1723858470
transform 1 0 2277 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_31
timestamp 1723858470
transform 1 0 1653 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_32
timestamp 1723858470
transform 1 0 3279 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_33
timestamp 1723858470
transform 1 0 3743 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_34
timestamp 1723858470
transform 1 0 3147 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_35
timestamp 1723858470
transform 1 0 2683 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_36
timestamp 1723858470
transform 1 0 2031 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_37
timestamp 1723858470
transform 1 0 2495 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_38
timestamp 1723858470
transform 1 0 1899 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_39
timestamp 1723858470
transform 1 0 1435 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_40
timestamp 1723858470
transform 1 0 5775 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_41
timestamp 1723858470
transform 1 0 6239 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_42
timestamp 1723858470
transform 1 0 5643 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_43
timestamp 1723858470
transform 1 0 5179 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_44
timestamp 1723858470
transform 1 0 4527 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_45
timestamp 1723858470
transform 1 0 4991 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_46
timestamp 1723858470
transform 1 0 4395 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_47
timestamp 1723858470
transform 1 0 3931 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_48
timestamp 1723858470
transform 1 0 18255 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_49
timestamp 1723858470
transform 1 0 18719 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_50
timestamp 1723858470
transform 1 0 18123 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_51
timestamp 1723858470
transform 1 0 17659 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_52
timestamp 1723858470
transform 1 0 17007 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_53
timestamp 1723858470
transform 1 0 17471 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_54
timestamp 1723858470
transform 1 0 16875 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_55
timestamp 1723858470
transform 1 0 16411 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_56
timestamp 1723858470
transform 1 0 20997 0 1 1233
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_57
timestamp 1723858470
transform 1 0 20373 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_58
timestamp 1723858470
transform 1 0 19749 0 1 985
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_59
timestamp 1723858470
transform 1 0 19125 0 1 861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_60
timestamp 1723858470
transform 1 0 18501 0 1 737
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_61
timestamp 1723858470
transform 1 0 17877 0 1 613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_62
timestamp 1723858470
transform 1 0 17253 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_63
timestamp 1723858470
transform 1 0 16629 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_64
timestamp 1723858470
transform 1 0 20751 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_65
timestamp 1723858470
transform 1 0 21215 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_66
timestamp 1723858470
transform 1 0 20619 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_67
timestamp 1723858470
transform 1 0 20155 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_68
timestamp 1723858470
transform 1 0 19503 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_69
timestamp 1723858470
transform 1 0 19967 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_70
timestamp 1723858470
transform 1 0 19371 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_71
timestamp 1723858470
transform 1 0 18907 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_72
timestamp 1723858470
transform 1 0 13509 0 1 737
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_73
timestamp 1723858470
transform 1 0 12885 0 1 613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_74
timestamp 1723858470
transform 1 0 12261 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_75
timestamp 1723858470
transform 1 0 11637 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_76
timestamp 1723858470
transform 1 0 15759 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_77
timestamp 1723858470
transform 1 0 16223 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_78
timestamp 1723858470
transform 1 0 15627 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_79
timestamp 1723858470
transform 1 0 15163 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_80
timestamp 1723858470
transform 1 0 14511 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_81
timestamp 1723858470
transform 1 0 14975 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_82
timestamp 1723858470
transform 1 0 14379 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_83
timestamp 1723858470
transform 1 0 13915 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_84
timestamp 1723858470
transform 1 0 13263 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_85
timestamp 1723858470
transform 1 0 13727 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_86
timestamp 1723858470
transform 1 0 13131 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_87
timestamp 1723858470
transform 1 0 12667 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_88
timestamp 1723858470
transform 1 0 12015 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_89
timestamp 1723858470
transform 1 0 12479 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_90
timestamp 1723858470
transform 1 0 11883 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_91
timestamp 1723858470
transform 1 0 11419 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_92
timestamp 1723858470
transform 1 0 16005 0 1 1233
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_93
timestamp 1723858470
transform 1 0 15381 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_94
timestamp 1723858470
transform 1 0 14757 0 1 985
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_95
timestamp 1723858470
transform 1 0 14133 0 1 861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_96
timestamp 1723858470
transform 1 0 30735 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_97
timestamp 1723858470
transform 1 0 31199 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_98
timestamp 1723858470
transform 1 0 30603 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_99
timestamp 1723858470
transform 1 0 30139 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_100
timestamp 1723858470
transform 1 0 29487 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_101
timestamp 1723858470
transform 1 0 29951 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_102
timestamp 1723858470
transform 1 0 29355 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_103
timestamp 1723858470
transform 1 0 28891 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_104
timestamp 1723858470
transform 1 0 28239 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_105
timestamp 1723858470
transform 1 0 28703 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_106
timestamp 1723858470
transform 1 0 28107 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_107
timestamp 1723858470
transform 1 0 27643 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_108
timestamp 1723858470
transform 1 0 26991 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_109
timestamp 1723858470
transform 1 0 27455 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_110
timestamp 1723858470
transform 1 0 26859 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_111
timestamp 1723858470
transform 1 0 26395 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_112
timestamp 1723858470
transform 1 0 28485 0 1 737
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_113
timestamp 1723858470
transform 1 0 27861 0 1 613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_114
timestamp 1723858470
transform 1 0 27237 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_115
timestamp 1723858470
transform 1 0 26613 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_116
timestamp 1723858470
transform 1 0 30981 0 1 1233
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_117
timestamp 1723858470
transform 1 0 30357 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_118
timestamp 1723858470
transform 1 0 29733 0 1 985
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_119
timestamp 1723858470
transform 1 0 29109 0 1 861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_120
timestamp 1723858470
transform 1 0 25989 0 1 1233
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_121
timestamp 1723858470
transform 1 0 25365 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_122
timestamp 1723858470
transform 1 0 24741 0 1 985
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_123
timestamp 1723858470
transform 1 0 24117 0 1 861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_124
timestamp 1723858470
transform 1 0 23493 0 1 737
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_125
timestamp 1723858470
transform 1 0 22869 0 1 613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_126
timestamp 1723858470
transform 1 0 22245 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_127
timestamp 1723858470
transform 1 0 21621 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_128
timestamp 1723858470
transform 1 0 23247 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_129
timestamp 1723858470
transform 1 0 23711 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_130
timestamp 1723858470
transform 1 0 23115 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_131
timestamp 1723858470
transform 1 0 22651 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_132
timestamp 1723858470
transform 1 0 21999 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_133
timestamp 1723858470
transform 1 0 22463 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_134
timestamp 1723858470
transform 1 0 21867 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_135
timestamp 1723858470
transform 1 0 21403 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_136
timestamp 1723858470
transform 1 0 25743 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_137
timestamp 1723858470
transform 1 0 26207 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_138
timestamp 1723858470
transform 1 0 25611 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_139
timestamp 1723858470
transform 1 0 25147 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_140
timestamp 1723858470
transform 1 0 24495 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_141
timestamp 1723858470
transform 1 0 24959 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_142
timestamp 1723858470
transform 1 0 24363 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_143
timestamp 1723858470
transform 1 0 23899 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_144
timestamp 1723858470
transform 1 0 40719 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_145
timestamp 1723858470
transform 1 0 41183 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_146
timestamp 1723858470
transform 1 0 40587 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_147
timestamp 1723858470
transform 1 0 40123 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_148
timestamp 1723858470
transform 1 0 39471 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_149
timestamp 1723858470
transform 1 0 39935 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_150
timestamp 1723858470
transform 1 0 39339 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_151
timestamp 1723858470
transform 1 0 38875 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_152
timestamp 1723858470
transform 1 0 38223 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_153
timestamp 1723858470
transform 1 0 38687 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_154
timestamp 1723858470
transform 1 0 38091 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_155
timestamp 1723858470
transform 1 0 37627 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_156
timestamp 1723858470
transform 1 0 36975 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_157
timestamp 1723858470
transform 1 0 37439 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_158
timestamp 1723858470
transform 1 0 36843 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_159
timestamp 1723858470
transform 1 0 36379 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_160
timestamp 1723858470
transform 1 0 40965 0 1 1233
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_161
timestamp 1723858470
transform 1 0 40341 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_162
timestamp 1723858470
transform 1 0 39717 0 1 985
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_163
timestamp 1723858470
transform 1 0 39093 0 1 861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_164
timestamp 1723858470
transform 1 0 38469 0 1 737
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_165
timestamp 1723858470
transform 1 0 37845 0 1 613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_166
timestamp 1723858470
transform 1 0 37221 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_167
timestamp 1723858470
transform 1 0 36597 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_168
timestamp 1723858470
transform 1 0 35727 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_169
timestamp 1723858470
transform 1 0 36191 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_170
timestamp 1723858470
transform 1 0 35595 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_171
timestamp 1723858470
transform 1 0 35131 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_172
timestamp 1723858470
transform 1 0 34479 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_173
timestamp 1723858470
transform 1 0 34943 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_174
timestamp 1723858470
transform 1 0 34347 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_175
timestamp 1723858470
transform 1 0 33883 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_176
timestamp 1723858470
transform 1 0 33231 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_177
timestamp 1723858470
transform 1 0 33695 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_178
timestamp 1723858470
transform 1 0 33099 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_179
timestamp 1723858470
transform 1 0 32635 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_180
timestamp 1723858470
transform 1 0 31983 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_181
timestamp 1723858470
transform 1 0 32447 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_182
timestamp 1723858470
transform 1 0 31851 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_183
timestamp 1723858470
transform 1 0 31387 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_184
timestamp 1723858470
transform 1 0 35973 0 1 1233
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_185
timestamp 1723858470
transform 1 0 35349 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_186
timestamp 1723858470
transform 1 0 34725 0 1 985
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_187
timestamp 1723858470
transform 1 0 34101 0 1 861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_188
timestamp 1723858470
transform 1 0 33477 0 1 737
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_189
timestamp 1723858470
transform 1 0 32853 0 1 613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_190
timestamp 1723858470
transform 1 0 32229 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_27_191
timestamp 1723858470
transform 1 0 31605 0 1 365
box 0 0 1 1
<< labels >>
rlabel metal3 s 0 372 41310 432 4 sel_0
port 1 nsew
rlabel metal3 s 0 496 41310 556 4 sel_1
port 2 nsew
rlabel metal3 s 0 620 41310 680 4 sel_2
port 3 nsew
rlabel metal3 s 0 744 41310 804 4 sel_3
port 4 nsew
rlabel metal3 s 0 868 41310 928 4 sel_4
port 5 nsew
rlabel metal3 s 0 992 41310 1052 4 sel_5
port 6 nsew
rlabel metal3 s 0 1116 41310 1176 4 sel_6
port 7 nsew
rlabel metal3 s 0 1240 41310 1300 4 sel_7
port 8 nsew
rlabel metal3 s 14429 1978 14527 2076 4 gnd
port 9 nsew
rlabel metal3 s 14478 2027 14478 2027 4 gnd
rlabel metal3 s 10685 1978 10783 2076 4 gnd
port 9 nsew
rlabel metal3 s 16925 1978 17023 2076 4 gnd
port 9 nsew
rlabel metal3 s 6941 1978 7039 2076 4 gnd
port 9 nsew
rlabel metal3 s 19421 1978 19519 2076 4 gnd
port 9 nsew
rlabel metal3 s 5693 1978 5791 2076 4 gnd
port 9 nsew
rlabel metal3 s 5742 2027 5742 2027 4 gnd
rlabel metal3 s 18173 1978 18271 2076 4 gnd
port 9 nsew
rlabel metal3 s 18222 2027 18222 2027 4 gnd
rlabel metal3 s 26909 1978 27007 2076 4 gnd
port 9 nsew
rlabel metal3 s 26958 2027 26958 2027 4 gnd
rlabel metal3 s 34397 1978 34495 2076 4 gnd
port 9 nsew
rlabel metal3 s 34446 2027 34446 2027 4 gnd
rlabel metal3 s 9437 1978 9535 2076 4 gnd
port 9 nsew
rlabel metal3 s 11933 1978 12031 2076 4 gnd
port 9 nsew
rlabel metal3 s 25661 1978 25759 2076 4 gnd
port 9 nsew
rlabel metal3 s 30653 1978 30751 2076 4 gnd
port 9 nsew
rlabel metal3 s 30702 2027 30702 2027 4 gnd
rlabel metal3 s 29405 1978 29503 2076 4 gnd
port 9 nsew
rlabel metal3 s 33149 1978 33247 2076 4 gnd
port 9 nsew
rlabel metal3 s 38141 1978 38239 2076 4 gnd
port 9 nsew
rlabel metal3 s 38190 2027 38190 2027 4 gnd
rlabel metal3 s 3197 1978 3295 2076 4 gnd
port 9 nsew
rlabel metal3 s 3246 2027 3246 2027 4 gnd
rlabel metal3 s 1949 1978 2047 2076 4 gnd
port 9 nsew
rlabel metal3 s 1998 2027 1998 2027 4 gnd
rlabel metal3 s 21917 1978 22015 2076 4 gnd
port 9 nsew
rlabel metal3 s 23165 1978 23263 2076 4 gnd
port 9 nsew
rlabel metal3 s 31901 1978 31999 2076 4 gnd
port 9 nsew
rlabel metal3 s 13181 1978 13279 2076 4 gnd
port 9 nsew
rlabel metal3 s 40637 1978 40735 2076 4 gnd
port 9 nsew
rlabel metal3 s 8189 1978 8287 2076 4 gnd
port 9 nsew
rlabel metal3 s 39389 1978 39487 2076 4 gnd
port 9 nsew
rlabel metal3 s 4445 1978 4543 2076 4 gnd
port 9 nsew
rlabel metal3 s 4494 2027 4494 2027 4 gnd
rlabel metal3 s 15677 1978 15775 2076 4 gnd
port 9 nsew
rlabel metal3 s 35645 1978 35743 2076 4 gnd
port 9 nsew
rlabel metal3 s 36893 1978 36991 2076 4 gnd
port 9 nsew
rlabel metal3 s 20669 1978 20767 2076 4 gnd
port 9 nsew
rlabel metal3 s 20718 2027 20718 2027 4 gnd
rlabel metal3 s 24413 1978 24511 2076 4 gnd
port 9 nsew
rlabel metal3 s 24462 2027 24462 2027 4 gnd
rlabel metal3 s 28157 1978 28255 2076 4 gnd
port 9 nsew
rlabel metal3 s 10734 2027 10734 2027 4 gnd
rlabel metal1 s 21422 248 21450 1364 4 bl_out_4
port 10 nsew
rlabel metal1 s 26414 248 26442 1364 4 bl_out_5
port 11 nsew
rlabel metal1 s 31406 248 31434 1364 4 bl_out_6
port 12 nsew
rlabel metal1 s 36398 248 36426 1364 4 bl_out_7
port 13 nsew
rlabel metal1 s 21422 2624 21450 2680 4 bl_32
port 14 nsew
rlabel metal1 s 21886 2624 21914 2680 4 br_32
port 15 nsew
rlabel metal1 s 22482 2624 22510 2680 4 bl_33
port 16 nsew
rlabel metal1 s 22018 2624 22046 2680 4 br_33
port 17 nsew
rlabel metal1 s 22670 2624 22698 2680 4 bl_34
port 18 nsew
rlabel metal1 s 23134 2624 23162 2680 4 br_34
port 19 nsew
rlabel metal1 s 23730 2624 23758 2680 4 bl_35
port 20 nsew
rlabel metal1 s 23266 2624 23294 2680 4 br_35
port 21 nsew
rlabel metal1 s 23918 2624 23946 2680 4 bl_36
port 22 nsew
rlabel metal1 s 24382 2624 24410 2680 4 br_36
port 23 nsew
rlabel metal1 s 24978 2624 25006 2680 4 bl_37
port 24 nsew
rlabel metal1 s 24514 2624 24542 2680 4 br_37
port 25 nsew
rlabel metal1 s 25166 2624 25194 2680 4 bl_38
port 26 nsew
rlabel metal1 s 25630 2624 25658 2680 4 br_38
port 27 nsew
rlabel metal1 s 26226 2624 26254 2680 4 bl_39
port 28 nsew
rlabel metal1 s 25762 2624 25790 2680 4 br_39
port 29 nsew
rlabel metal1 s 26414 2624 26442 2680 4 bl_40
port 30 nsew
rlabel metal1 s 26878 2624 26906 2680 4 br_40
port 31 nsew
rlabel metal1 s 27474 2624 27502 2680 4 bl_41
port 32 nsew
rlabel metal1 s 27010 2624 27038 2680 4 br_41
port 33 nsew
rlabel metal1 s 27662 2624 27690 2680 4 bl_42
port 34 nsew
rlabel metal1 s 28126 2624 28154 2680 4 br_42
port 35 nsew
rlabel metal1 s 28722 2624 28750 2680 4 bl_43
port 36 nsew
rlabel metal1 s 28258 2624 28286 2680 4 br_43
port 37 nsew
rlabel metal1 s 28910 2624 28938 2680 4 bl_44
port 38 nsew
rlabel metal1 s 29374 2624 29402 2680 4 br_44
port 39 nsew
rlabel metal1 s 29970 2624 29998 2680 4 bl_45
port 40 nsew
rlabel metal1 s 29506 2624 29534 2680 4 br_45
port 41 nsew
rlabel metal1 s 30158 2624 30186 2680 4 bl_46
port 42 nsew
rlabel metal1 s 30622 2624 30650 2680 4 br_46
port 43 nsew
rlabel metal1 s 31218 2624 31246 2680 4 bl_47
port 44 nsew
rlabel metal1 s 30754 2624 30782 2680 4 br_47
port 45 nsew
rlabel metal1 s 31406 2624 31434 2680 4 bl_48
port 46 nsew
rlabel metal1 s 31870 2624 31898 2680 4 br_48
port 47 nsew
rlabel metal1 s 32466 2624 32494 2680 4 bl_49
port 48 nsew
rlabel metal1 s 32002 2624 32030 2680 4 br_49
port 49 nsew
rlabel metal1 s 32654 2624 32682 2680 4 bl_50
port 50 nsew
rlabel metal1 s 33118 2624 33146 2680 4 br_50
port 51 nsew
rlabel metal1 s 33714 2624 33742 2680 4 bl_51
port 52 nsew
rlabel metal1 s 33250 2624 33278 2680 4 br_51
port 53 nsew
rlabel metal1 s 33902 2624 33930 2680 4 bl_52
port 54 nsew
rlabel metal1 s 34366 2624 34394 2680 4 br_52
port 55 nsew
rlabel metal1 s 34962 2624 34990 2680 4 bl_53
port 56 nsew
rlabel metal1 s 34498 2624 34526 2680 4 br_53
port 57 nsew
rlabel metal1 s 35150 2624 35178 2680 4 bl_54
port 58 nsew
rlabel metal1 s 35614 2624 35642 2680 4 br_54
port 59 nsew
rlabel metal1 s 36210 2624 36238 2680 4 bl_55
port 60 nsew
rlabel metal1 s 35746 2624 35774 2680 4 br_55
port 61 nsew
rlabel metal1 s 36398 2624 36426 2680 4 bl_56
port 62 nsew
rlabel metal1 s 36862 2624 36890 2680 4 br_56
port 63 nsew
rlabel metal1 s 37458 2624 37486 2680 4 bl_57
port 64 nsew
rlabel metal1 s 36994 2624 37022 2680 4 br_57
port 65 nsew
rlabel metal1 s 37646 2624 37674 2680 4 bl_58
port 66 nsew
rlabel metal1 s 38110 2624 38138 2680 4 br_58
port 67 nsew
rlabel metal1 s 38706 2624 38734 2680 4 bl_59
port 68 nsew
rlabel metal1 s 38242 2624 38270 2680 4 br_59
port 69 nsew
rlabel metal1 s 38894 2624 38922 2680 4 bl_60
port 70 nsew
rlabel metal1 s 39358 2624 39386 2680 4 br_60
port 71 nsew
rlabel metal1 s 39954 2624 39982 2680 4 bl_61
port 72 nsew
rlabel metal1 s 39490 2624 39518 2680 4 br_61
port 73 nsew
rlabel metal1 s 40142 2624 40170 2680 4 bl_62
port 74 nsew
rlabel metal1 s 40606 2624 40634 2680 4 br_62
port 75 nsew
rlabel metal1 s 41202 2624 41230 2680 4 bl_63
port 76 nsew
rlabel metal1 s 40738 2624 40766 2680 4 br_63
port 77 nsew
rlabel metal1 s 20174 2624 20202 2680 4 bl_30
port 78 nsew
rlabel metal1 s 20638 2624 20666 2680 4 br_30
port 79 nsew
rlabel metal1 s 21234 2624 21262 2680 4 bl_31
port 80 nsew
rlabel metal1 s 20770 2624 20798 2680 4 br_31
port 81 nsew
rlabel metal1 s 1454 248 1482 1364 4 bl_out_0
port 82 nsew
rlabel metal1 s 6446 248 6474 1364 4 bl_out_1
port 83 nsew
rlabel metal1 s 11438 248 11466 1364 4 bl_out_2
port 84 nsew
rlabel metal1 s 16430 248 16458 1364 4 bl_out_3
port 85 nsew
rlabel metal1 s 1454 2624 1482 2680 4 bl_0
port 86 nsew
rlabel metal1 s 1918 2624 1946 2680 4 br_0
port 87 nsew
rlabel metal1 s 2514 2624 2542 2680 4 bl_1
port 88 nsew
rlabel metal1 s 2050 2624 2078 2680 4 br_1
port 89 nsew
rlabel metal1 s 2702 2624 2730 2680 4 bl_2
port 90 nsew
rlabel metal1 s 3166 2624 3194 2680 4 br_2
port 91 nsew
rlabel metal1 s 3762 2624 3790 2680 4 bl_3
port 92 nsew
rlabel metal1 s 3298 2624 3326 2680 4 br_3
port 93 nsew
rlabel metal1 s 3950 2624 3978 2680 4 bl_4
port 94 nsew
rlabel metal1 s 4414 2624 4442 2680 4 br_4
port 95 nsew
rlabel metal1 s 5010 2624 5038 2680 4 bl_5
port 96 nsew
rlabel metal1 s 4546 2624 4574 2680 4 br_5
port 97 nsew
rlabel metal1 s 5198 2624 5226 2680 4 bl_6
port 98 nsew
rlabel metal1 s 5662 2624 5690 2680 4 br_6
port 99 nsew
rlabel metal1 s 6258 2624 6286 2680 4 bl_7
port 100 nsew
rlabel metal1 s 5794 2624 5822 2680 4 br_7
port 101 nsew
rlabel metal1 s 6446 2624 6474 2680 4 bl_8
port 102 nsew
rlabel metal1 s 6910 2624 6938 2680 4 br_8
port 103 nsew
rlabel metal1 s 7506 2624 7534 2680 4 bl_9
port 104 nsew
rlabel metal1 s 7042 2624 7070 2680 4 br_9
port 105 nsew
rlabel metal1 s 7694 2624 7722 2680 4 bl_10
port 106 nsew
rlabel metal1 s 8158 2624 8186 2680 4 br_10
port 107 nsew
rlabel metal1 s 8754 2624 8782 2680 4 bl_11
port 108 nsew
rlabel metal1 s 8290 2624 8318 2680 4 br_11
port 109 nsew
rlabel metal1 s 8942 2624 8970 2680 4 bl_12
port 110 nsew
rlabel metal1 s 9406 2624 9434 2680 4 br_12
port 111 nsew
rlabel metal1 s 10002 2624 10030 2680 4 bl_13
port 112 nsew
rlabel metal1 s 9538 2624 9566 2680 4 br_13
port 113 nsew
rlabel metal1 s 10190 2624 10218 2680 4 bl_14
port 114 nsew
rlabel metal1 s 10654 2624 10682 2680 4 br_14
port 115 nsew
rlabel metal1 s 11250 2624 11278 2680 4 bl_15
port 116 nsew
rlabel metal1 s 10786 2624 10814 2680 4 br_15
port 117 nsew
rlabel metal1 s 11438 2624 11466 2680 4 bl_16
port 118 nsew
rlabel metal1 s 11902 2624 11930 2680 4 br_16
port 119 nsew
rlabel metal1 s 12498 2624 12526 2680 4 bl_17
port 120 nsew
rlabel metal1 s 12034 2624 12062 2680 4 br_17
port 121 nsew
rlabel metal1 s 12686 2624 12714 2680 4 bl_18
port 122 nsew
rlabel metal1 s 13150 2624 13178 2680 4 br_18
port 123 nsew
rlabel metal1 s 13746 2624 13774 2680 4 bl_19
port 124 nsew
rlabel metal1 s 13282 2624 13310 2680 4 br_19
port 125 nsew
rlabel metal1 s 13934 2624 13962 2680 4 bl_20
port 126 nsew
rlabel metal1 s 14398 2624 14426 2680 4 br_20
port 127 nsew
rlabel metal1 s 14994 2624 15022 2680 4 bl_21
port 128 nsew
rlabel metal1 s 14530 2624 14558 2680 4 br_21
port 129 nsew
rlabel metal1 s 15182 2624 15210 2680 4 bl_22
port 130 nsew
rlabel metal1 s 15646 2624 15674 2680 4 br_22
port 131 nsew
rlabel metal1 s 16242 2624 16270 2680 4 bl_23
port 132 nsew
rlabel metal1 s 15778 2624 15806 2680 4 br_23
port 133 nsew
rlabel metal1 s 16430 2624 16458 2680 4 bl_24
port 134 nsew
rlabel metal1 s 16894 2624 16922 2680 4 br_24
port 135 nsew
rlabel metal1 s 17490 2624 17518 2680 4 bl_25
port 136 nsew
rlabel metal1 s 17026 2624 17054 2680 4 br_25
port 137 nsew
rlabel metal1 s 17678 2624 17706 2680 4 bl_26
port 138 nsew
rlabel metal1 s 18142 2624 18170 2680 4 br_26
port 139 nsew
rlabel metal1 s 18738 2624 18766 2680 4 bl_27
port 140 nsew
rlabel metal1 s 18274 2624 18302 2680 4 br_27
port 141 nsew
rlabel metal1 s 18926 2624 18954 2680 4 bl_28
port 142 nsew
rlabel metal1 s 19390 2624 19418 2680 4 br_28
port 143 nsew
rlabel metal1 s 19986 2624 20014 2680 4 bl_29
port 144 nsew
rlabel metal1 s 19522 2624 19550 2680 4 br_29
port 145 nsew
rlabel metal1 s 1918 124 1946 1364 4 br_out_0
port 146 nsew
rlabel metal1 s 11902 124 11930 1364 4 br_out_2
port 147 nsew
rlabel metal1 s 6910 124 6938 1364 4 br_out_1
port 148 nsew
rlabel metal1 s 16894 124 16922 1364 4 br_out_3
port 149 nsew
rlabel metal1 s 21886 124 21914 1364 4 br_out_4
port 150 nsew
rlabel metal1 s 31870 124 31898 1364 4 br_out_6
port 151 nsew
rlabel metal1 s 26878 124 26906 1364 4 br_out_5
port 152 nsew
rlabel metal1 s 36862 124 36890 1364 4 br_out_7
port 153 nsew
<< properties >>
string FIXED_BBOX 40719 87 40785 161
string GDS_END 1048072
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 941686
<< end >>

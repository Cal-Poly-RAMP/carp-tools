magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -36 679 2672 1471
<< pwell >>
rect 2500 25 2602 159
<< psubdiff >>
rect 2526 109 2576 133
rect 2526 75 2534 109
rect 2568 75 2576 109
rect 2526 51 2576 75
<< nsubdiff >>
rect 2526 1339 2576 1363
rect 2526 1305 2534 1339
rect 2568 1305 2576 1339
rect 2526 1281 2576 1305
<< psubdiffcont >>
rect 2534 75 2568 109
<< nsubdiffcont >>
rect 2534 1305 2568 1339
<< poly >>
rect 114 740 144 907
rect 48 724 144 740
rect 48 690 64 724
rect 98 690 144 724
rect 48 674 144 690
rect 114 507 144 674
<< polycont >>
rect 64 690 98 724
<< locali >>
rect 0 1397 2636 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 490 1130 524 1397
rect 706 1130 740 1397
rect 922 1130 956 1397
rect 1138 1130 1172 1397
rect 1354 1130 1388 1397
rect 1570 1130 1604 1397
rect 1786 1130 1820 1397
rect 2002 1130 2036 1397
rect 2218 1130 2252 1397
rect 2430 1130 2464 1397
rect 2534 1339 2568 1397
rect 2534 1289 2568 1305
rect 64 724 98 740
rect 64 674 98 690
rect 1246 724 1280 1096
rect 1246 690 1297 724
rect 1246 318 1280 690
rect 62 17 96 218
rect 274 17 308 218
rect 490 17 524 218
rect 706 17 740 218
rect 922 17 956 218
rect 1138 17 1172 218
rect 1354 17 1388 218
rect 1570 17 1604 218
rect 1786 17 1820 218
rect 2002 17 2036 218
rect 2218 17 2252 218
rect 2430 17 2464 218
rect 2534 109 2568 125
rect 2534 17 2568 75
rect 0 -17 2636 17
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_16  sky130_sram_2kbyte_1rw1r_32x512_8_contact_16_0
timestamp 1723858470
transform 1 0 48 0 1 674
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_28  sky130_sram_2kbyte_1rw1r_32x512_8_contact_28_0
timestamp 1723858470
transform 1 0 2526 0 1 1281
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_29  sky130_sram_2kbyte_1rw1r_32x512_8_contact_29_0
timestamp 1723858470
transform 1 0 2526 0 1 51
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m22_w2_000_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m22_w2_000_sli_dli_da_p_0
timestamp 1723858470
transform 1 0 54 0 1 51
box -26 -26 2444 456
use sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m22_w2_000_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m22_w2_000_sli_dli_da_p_0
timestamp 1723858470
transform 1 0 54 0 1 963
box -59 -56 2477 454
<< labels >>
rlabel locali s 81 707 81 707 4 A
rlabel locali s 1280 707 1280 707 4 Z
rlabel locali s 1318 0 1318 0 4 gnd
rlabel locali s 1318 1414 1318 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 2636 1414
string GDS_END 106162
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 102884
<< end >>
